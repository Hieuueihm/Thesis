module ci_top #(
    parameter ROWS = 30,
    parameter COLS = 30
) (
    input clk,
    input rst_n,
    input [7:0] grayscale_i,
    input i_valid,
    output [15:0] r2_bit_one_o,
    output [15:0] r2_bit_zero_o,
    output done_r2,
    output [15:0] r4_bit_one_o,
    output [15:0] r4_bit_zero_o,
    output done_r4,
    output [15:0] r6_bit_one_o,
    output [15:0] r6_bit_zero_o,
    output done_r6,
    output [15:0] R8_bit_one_o,
    output [15:0] R8_bit_zero_o,
    output done_R8
);


  wire [7:0] d0_o, d1_o, d2_o, d3_o, d4_o, d5_o, d6_o, d7_o, d8_o;
  wire prepare_;
  // preparation == buffer
  preparation #(
      .DEPTH(COLS)
  ) median_PREPARATION (
      .clk(clk),
      .rst_n(rst_n),
      .i_valid(i_valid),
      .data_i(grayscale_i),
      .data0_o(d0_o),
      .data1_o(d1_o),
      .data2_o(d2_o),
      .data3_o(d3_o),
      .data4_o(d4_o),
      .data5_o(d5_o),
      .data6_o(d6_o),
      .data7_o(d7_o),
      .data8_o(d8_o),
      .(prepare_)
  );
  // median = datamodulat + calc
  wire median_;
  wire [7:0] median_o;
  median_filter_3x3 #(
      .ROWS(ROWS),
      .COLS(COLS)
  ) median_FILTER_3x3 (
      .clk(clk),
      .rst_n(rst_n),
      .i_valid(prepare_),
      .d0_i(d0_o),
      .d1_i(d1_o),
      .d2_i(d2_o),
      .d3_i(d3_o),
      .d4_i(d4_o),
      .d5_i(d5_o),
      .d6_i(d6_o),
      .d7_i(d7_o),
      .d8_i(d8_o),
      .median_o(median_o),
      .(median_)
  );
  // buffer 16 rows;
  wire [7:0] data0_o;
  wire [7:0] data1_o;
  wire [7:0] data2_o;
  wire [7:0] data3_o;
  wire [7:0] data4_o;
  wire [7:0] data5_o;
  wire [7:0] data6_o;
  wire [7:0] data7_o;
  wire [7:0] data8_o;
  wire [7:0] data9_o, data10_o, data11_o, data12_o, data13_o, data14_o, data15_o, data16_o;
  wire buffer_16_;
  buffer_16_rows #(
      .DEPTH(COLS)
  ) BUFFER_16_ROWS (
      .clk(clk),
      .rst_n(rst_n),
      .i_valid(median_),
      .data_i(median_o),
      .data0_o(data0_o),
      .data1_o(data1_o),
      .data2_o(data2_o),
      .data3_o(data3_o),
      .data4_o(data4_o),
      .data5_o(data5_o),
      .data6_o(data6_o),
      .data7_o(data7_o),
      .data8_o(data8_o),
      .data9_o(data9_o),
      .data10_o(data10_o),
      .data11_o(data11_o),
      .data12_o(data12_o),
      .data13_o(data13_o),
      .data14_o(data14_o),
      .data15_o(data15_o),
      .data16_o(data16_o),
      .(buffer_16_)
  );



  // // ci calculation
  // r2_top #(.COLS(COLS),
  // .ROWS(ROWS))
  // r2_TOP
  // (
  // .clk(clk),
  // .rst_n(rst_n),
  // .i_valid(buffer_16_),
  // .S1(data12_o),
  // .S2(data13_o),
  // .S3(data14_o),
  // .S4(data15_o),
  // .S5(data16_o),
  // .(done_r2),
  // .bit_one_o(r2_bit_one_o),
  // .bit_zero_o(r2_bit_zero_o));

  // r4_top #(.COLS(COLS),
  // .ROWS(ROWS))
  // r4_TOP
  // (
  // .clk(clk),
  // .rst_n(rst_n),
  // .i_valid(buffer_16_),
  // .S1(data8_o),
  // .S2(data9_o),
  // .S3(data10_o),
  // .S4(data11_o),
  // .S5(data12_o),
  // .S6(data13_o),
  // .S7(data14_o),
  // .S8(data15_o),
  // .S9(data16_o),
  // .(done_r4),
  // .bit_one_o(r4_bit_one_o),
  // .bit_zero_o(r4_bit_zero_o));

  // r6_top #(.COLS(COLS),
  // .ROWS(ROWS))
  // r6_TOP
  // (
  // .clk(clk),
  // .rst_n(rst_n),
  // .i_valid(buffer_16_),
  // .S1(data4_o),
  // .S2(data5_o),
  // .S3(data6_o),
  // .S4(data7_o),
  // .S5(data8_o),
  // .S6(data9_o),
  // .S7(data10_o),
  // .S8(data11_o),
  // .S9(data12_o),
  // .S10(data13_o),
  // .S11(data14_o),
  // .S12(data15_o),
  // .S13(data16_o),
  // .(done_r6),
  // .bit_one_o(r6_bit_one_o),
  // .bit_zero_o(r6_bit_zero_o));

  // R8_top #(.COLS(COLS),
  // .ROWS(ROWS))
  // R8_TOP
  // (
  // .clk(clk),
  // .rst_n(rst_n),
  // .i_valid(buffer_16_),
  // .S1(data0_o),
  // .S2(data1_o),
  // .S3(data2_o),
  // .S4(data3_o),
  // .S5(data4_o),
  // .S6(data5_o),
  // .S7(data6_o),
  // .S8(data7_o),
  // .S9(data8_o),
  // .S10(data9_o),
  // .S11(data10_o),
  // .S12(data11_o),
  // .S13(data12_o),
  // .S14(data13_o),
  // .S15(data14_o),
  // .S16(data15_o),
  // .S17(data16_o),
  // .(done_R8),
  // .bit_one_o(R8_bit_one_o),
  // .bit_zero_o(R8_bit_zero_o));


endmodule
