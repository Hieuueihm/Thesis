module window_buffer_7x7 (
    input clk,
    input rst_n,
    input data_valid_i,
    input start_i,
    input [7:0] S1_i,
    S2_i,
    S3_i,
    S4_i,
    S5_i,
    S6_i,
    S7_i,
    input [8:0] IMG_SIZE_I,
    output [7:0] S1_o,
    S2_o,
    S3_o,
    S4_o,
    S5_o,
    S6_o,
    S7_o,
    S8_o,
    S9_o,
    S10_o,
    S11_o,
    S12_o,
    S13_o,
    S14_o,
    S15_o,
    S16_o,
    S17_o,
    S18_o,
    S19_o,
    S20_o,
    S21_o,
    S22_o,
    S23_o,
    S24_o,
    S25_o,
    S26_o,
    S27_o,
    S28_o,
    S29_o,
    S30_o,
    S31_o,
    S32_o,
    S33_o,
    S34_o,
    S35_o,
    S36_o,
    S37_o,
    S38_o,
    S39_o,
    S40_o,
    S41_o,
    S42_o,
    S43_o,
    S44_o,
    S45_o,
    S46_o,
    S47_o,
    S48_o,
    S49_o,
    output data_valid_o,
    output finish_o
);
  wire i_row_eq_max, i_col_eq_max, i_col_ge_threshold;
  wire count_en;
  wire reset_en;
  window_buffer_controller inst_window_buffer_controller_7x7 (
      .clk                (clk),
      .rst_n              (rst_n),
      .start_i       (start_i),
      .i_row_eq_max       (i_row_eq_max),
      .i_col_eq_max       (i_col_eq_max),
      .i_col_ge_threshold (i_col_ge_threshold),
      .count_en           (count_en),
      .finish_o           (finish_o),
      .data_valid_o       (data_valid_o),
      .reset_en           (reset_en)
    );


  window_buffer_7x7_datapath inst_window_buffer_7x7_datapath
    (
      .clk                (clk),
      .rst_n              (rst_n),
      .count_en           (count_en),
      .S1_i               (S1_i),
      .S2_i               (S2_i),
      .S3_i               (S3_i),
      .S4_i               (S4_i),
      .S5_i               (S5_i),
      .S6_i               (S6_i),
      .S7_i               (S7_i),
      .data_valid_i      (data_valid_i),
      .IMG_SIZE_I         (IMG_SIZE_I),
      .i_row_eq_max       (i_row_eq_max),
      .S1_o               (S1_o),
      .S2_o               (S2_o),
      .S3_o               (S3_o),
      .S4_o               (S4_o),
      .S5_o               (S5_o),
      .S6_o               (S6_o),
      .S7_o               (S7_o),
      .S8_o               (S8_o),
      .S9_o               (S9_o),
      .S10_o              (S10_o),
      .S11_o              (S11_o),
      .S12_o              (S12_o),
      .S13_o              (S13_o),
      .S14_o              (S14_o),
      .S15_o              (S15_o),
      .S16_o              (S16_o),
      .S17_o              (S17_o),
      .S18_o              (S18_o),
      .S19_o              (S19_o),
      .S20_o              (S20_o),
      .S21_o              (S21_o),
      .S22_o              (S22_o),
      .S23_o              (S23_o),
      .S24_o              (S24_o),
      .S25_o              (S25_o),
      .S26_o              (S26_o),
      .S27_o              (S27_o),
      .S28_o              (S28_o),
      .S29_o              (S29_o),
      .S30_o              (S30_o),
      .S31_o              (S31_o),
      .S32_o              (S32_o),
      .S33_o              (S33_o),
      .S34_o              (S34_o),
      .S35_o              (S35_o),
      .S36_o              (S36_o),
      .S37_o              (S37_o),
      .S38_o              (S38_o),
      .S39_o              (S39_o),
      .S40_o              (S40_o),
      .S41_o              (S41_o),
      .S42_o              (S42_o),
      .S43_o              (S43_o),
      .S44_o              (S44_o),
      .S45_o              (S45_o),
      .S46_o              (S46_o),
      .S47_o              (S47_o),
      .S48_o              (S48_o),
      .S49_o              (S49_o),
      .i_col_eq_max       (i_col_eq_max),
      .i_col_ge_threshold (i_col_ge_threshold),
      .reset_en           (reset_en)
    );


endmodule
