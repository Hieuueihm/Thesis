module Serialiser (input clk,
                   input rst,
                   input done_i,
                   input [9:0] i_col,
                   input [7:0] S1,
                   S2,
                   S3,
                   S4,
                   S5,
                   S6,
                   S7,
                   S8,
                   S9,
                   S10,
                   S11,
                   S12,
                   S13,
                   S14,
                   S15,
                   S16,
                   S17,
                   S18,
                   S19,
                   S20,
                   S21,
                   S22,
                   S23,
                   S24,
                   S25,
                   output [7:0] S1_o,
                   S2_o,
                   S3_o,
                   S4_o,
                   S5_o,
                   output done_o,
                   output [2:0] o_select_o);
    
    wire [2:0] o_select_tmp;
    assign o_select_o = o_select_tmp;
    Serialiser_controller CONTROLLER
    (
    .clk(clk),
    .rst(rst),
    .i_col(i_col),
    .done_i(done_i),
    .o_select(o_select_tmp),
    .done_o(done_o));
    Serialiser_datapath DATAPATH(
    .clk(clk),
    .rst(rst),
    .S1(S1),
    .S2(S2),
    .S3(S3),
    .S4(S4),
    .S5(S5),
    .S6(S6),
    .S7(S7),
    .S8(S8),
    .S9(S9),
    .S10(S10),
    .S11(S11),
    .S12(S12),
    .S13(S13),
    .S14(S14),
    .S15(S15),
    .S16(S16),
    .S17(S17),
    .S18(S18),
    .S19(S19),
    .S20(S20),
    .S21(S21),
    .S22(S22),
    .S23(S23),
    .S24(S24),
    .S25(S25),
    .o_select(o_select_tmp),
    .S1_o(S1_o),
    .S2_o(S2_o),
    .S3_o(S3_o),
    .S4_o(S4_o),
    .S5_o(S5_o));
    
    
endmodule
