module sum_cumulative_top (input clk,
                           input rst,
                           input done_i,
                           input [9:0] i_col,
                           input [7:0] S1,
                           S2,
                           S3,
                           S4,
                           S5,
                           S6,
                           S7,
                           S8,
                           S9,
                           S10,
                           S11,
                           S12,
                           S13,
                           S14,
                           S15,
                           S16,
                           S17,
                           S18,
                           S19,
                           S20,
                           S21,
                           S22,
                           S23,
                           S24,
                           S25,
                           output done_o,
                           output [12:0] sum_o);
    
    
    wire [7:0]  S1_o, S2_o, S3_o, S4_o, S5_o;
    wire  done_o_temp;
    wire [2:0] o_select_o_temp;
    
    Serialiser SERIALISER(
    .clk(clk),
    .rst(rst),
    .done_i(done_i),
    .i_col(i_col),
    .S1(S1),
    .S2(S2),
    .S3(S3),
    .S4(S4),
    .S5(S5),
    .S6(S6),
    .S7(S7),
    .S8(S8),
    .S9(S9),
    .S10(S10),
    .S11(S11),
    .S12(S12),
    .S13(S13),
    .S14(S14),
    .S15(S15),
    .S16(S16),
    .S17(S17),
    .S18(S18),
    .S19(S19),
    .S20(S20),
    .S21(S21),
    .S22(S22),
    .S23(S23),
    .S24(S24),
    .S25(S25),
    .S1_o(S1_o),
    .S2_o(S2_o),
    .S3_o(S3_o),
    .S4_o(S4_o),
    .S5_o(S5_o),
    .done_o(done_o_temp),
    .o_select_o(o_select_o_temp));
    
    sum_cumulative SUM(
    .clk(clk),
    .rst(rst),
    .done_i(done_o_temp),
    .o_select_i(o_select_o_temp),
    .S1(S1_o),
    .S2(S2_o),
    .S3(S3_o),
    .S4(S4_o),
    .S5(S5_o),
    .sum_o(sum_o),
    .done_o(done_o));
    
endmodule
