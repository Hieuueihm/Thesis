module Data_modulate_17x17 #(
    parameter ROWS,
    parameter COLS
) (
    input clk,
    input rst,
    input done_i,
    input [7:0] data0_i,
    data1_i,
    data2_i,
    data3_i,
    data4_i,
    data5_i,
    data6_i,
    data7_i,
    data8_i,
    data9_i,
    data10_i,
    data11_i,
    data12_i,
    data13_i,
    data14_i,
    data15_i,
    data16_i,
    output reg [7:0] data0_o,
    data1_o,
    data2_o,
    data3_o,
    data4_o,
    data5_o,
    data6_o,
    data7_o,
    data8_o,
    data9_o,
    data10_o,
    data11_o,
    data12_o,
    data13_o,
    data14_o,
    data15_o,
    data16_o,
    data17_o,
    data18_o,
    data19_o,
    data20_o,
    data21_o,
    data22_o,
    data23_o,
    data24_o,
    data25_o,
    data26_o,
    data27_o,
    data28_o,
    data29_o,
    data30_o,
    data31_o,
    data32_o,
    data33_o,
    data34_o,
    data35_o,
    data36_o,
    data37_o,
    data38_o,
    data39_o,
    data40_o,
    data41_o,
    data42_o,
    data43_o,
    data44_o,
    data45_o,
    data46_o,
    data47_o,
    data48_o,
    data49_o,
    data50_o,
    data51_o,
    data52_o,
    data53_o,
    data54_o,
    data55_o,
    data56_o,
    data57_o,
    data58_o,
    data59_o,
    data60_o,
    data61_o,
    data62_o,
    data63_o,
    data64_o,
    data65_o,
    data66_o,
    data67_o,
    data68_o,
    data69_o,
    data70_o,
    data71_o,
    data72_o,
    data73_o,
    data74_o,
    data75_o,
    data76_o,
    data77_o,
    data78_o,
    data79_o,
    data80_o,
    data81_o,
    data82_o,
    data83_o,
    data84_o,
    data85_o,
    data86_o,
    data87_o,
    data88_o,
    data89_o,
    data90_o,
    data91_o,
    data92_o,
    data93_o,
    data94_o,
    data95_o,
    data96_o,
    data97_o,
    data98_o,
    data99_o,
    data100_o,
    data101_o,
    data102_o,
    data103_o,
    data104_o,
    data105_o,
    data106_o,
    data107_o,
    data108_o,
    data109_o,
    data110_o,
    data111_o,
    data112_o,
    data113_o,
    data114_o,
    data115_o,
    data116_o,
    data117_o,
    data118_o,
    data119_o,
    data120_o,
    data121_o,
    data122_o,
    data123_o,
    data124_o,
    data125_o,
    data126_o,
    data127_o,
    data128_o,
    data129_o,
    data130_o,
    data131_o,
    data132_o,
    data133_o,
    data134_o,
    data135_o,
    data136_o,
    data137_o,
    data138_o,
    data139_o,
    data140_o,
    data141_o,
    data142_o,
    data143_o,
    data144_o,
    data145_o,
    data146_o,
    data147_o,
    data148_o,
    data149_o,
    data150_o,
    data151_o,
    data152_o,
    data153_o,
    data154_o,
    data155_o,
    data156_o,
    data157_o,
    data158_o,
    data159_o,
    data160_o,
    data161_o,
    data162_o,
    data163_o,
    data164_o,
    data165_o,
    data166_o,
    data167_o,
    data168_o,
    data169_o,
    data170_o,
    data171_o,
    data172_o,
    data173_o,
    data174_o,
    data175_o,
    data176_o,
    data177_o,
    data178_o,
    data179_o,
    data180_o,
    data181_o,
    data182_o,
    data183_o,
    data184_o,
    data185_o,
    data186_o,
    data187_o,
    data188_o,
    data189_o,
    data190_o,
    data191_o,
    data192_o,
    data193_o,
    data194_o,
    data195_o,
    data196_o,
    data197_o,
    data198_o,
    data199_o,
    data200_o,
    data201_o,
    data202_o,
    data203_o,
    data204_o,
    data205_o,
    data206_o,
    data207_o,
    data208_o,
    data209_o,
    data210_o,
    data211_o,
    data212_o,
    data213_o,
    data214_o,
    data215_o,
    data216_o,
    data217_o,
    data218_o,
    data219_o,
    data220_o,
    data221_o,
    data222_o,
    data223_o,
    data224_o,
    data225_o,
    data226_o,
    data227_o,
    data228_o,
    data229_o,
    data230_o,
    data231_o,
    data232_o,
    data233_o,
    data234_o,
    data235_o,
    data236_o,
    data237_o,
    data238_o,
    data239_o,
    data240_o,
    data241_o,
    data242_o,
    data243_o,
    data244_o,
    data245_o,
    data246_o,
    data247_o,
    data248_o,
    data249_o,
    data250_o,
    data251_o,
    data252_o,
    data253_o,
    data254_o,
    data255_o,
    data256_o,
    data257_o,
    data258_o,
    data259_o,
    data260_o,
    data261_o,
    data262_o,
    data263_o,
    data264_o,
    data265_o,
    data266_o,
    data267_o,
    data268_o,
    data269_o,
    data270_o,
    data271_o,
    data272_o,
    data273_o,
    data274_o,
    data275_o,
    data276_o,
    data277_o,
    data278_o,
    data279_o,
    data280_o,
    data281_o,
    data282_o,
    data283_o,
    data284_o,
    data285_o,
    data286_o,
    data287_o,
    data288_o,
    output reg done_o
);

  reg [9:0] i_row, i_col;

  reg [7:0] i_counter;

  reg [7:0]
      data0,
      data1,
      data2,
      data3,
      data4,
      data5,
      data6,
      data7,
      data8,
      data9,
      data10,
      data11,
      data12,
      data13,
      data14,
      data15,
      data16,
      data17,
      data18,
      data19,
      data20,
      data21,
      data22,
      data23,
      data24,
      data25,
      data26,
      data27,
      data28,
      data29,
      data30,
      data31,
      data32,
      data33,
      data34,
      data35,
      data36,
      data37,
      data38,
      data39,
      data40,
      data41,
      data42,
      data43,
      data44,
      data45,
      data46,
      data47,
      data48,
      data49,
      data50,
      data51,
      data52,
      data53,
      data54,
      data55,
      data56,
      data57,
      data58,
      data59,
      data60,
      data61,
      data62,
      data63,
      data64,
      data65,
      data66,
      data67,
      data68,
      data69,
      data70,
      data71,
      data72,
      data73,
      data74,
      data75,
      data76,
      data77,
      data78,
      data79,
      data80,
      data81,
      data82,
      data83,
      data84,
      data85,
      data86,
      data87,
      data88,
      data89,
      data90,
      data91,
      data92,
      data93,
      data94,
      data95,
      data96,
      data97,
      data98,
      data99,
      data100,
      data101,
      data102,
      data103,
      data104,
      data105,
      data106,
      data107,
      data108,
      data109,
      data110,
      data111,
      data112,
      data113,
      data114,
      data115,
      data116,
      data117,
      data118,
      data119,
      data120,
      data121,
      data122,
      data123,
      data124,
      data125,
      data126,
      data127,
      data128,
      data129,
      data130,
      data131,
      data132,
      data133,
      data134,
      data135,
      data136,
      data137,
      data138,
      data139,
      data140,
      data141,
      data142,
      data143,
      data144,
      data145,
      data146,
      data147,
      data148,
      data149,
      data150,
      data151,
      data152,
      data153,
      data154,
      data155,
      data156,
      data157,
      data158,
      data159,
      data160,
      data161,
      data162,
      data163,
      data164,
      data165,
      data166,
      data167,
      data168,
      data169,
      data170,
      data171,
      data172,
      data173,
      data174,
      data175,
      data176,
      data177,
      data178,
      data179,
      data180,
      data181,
      data182,
      data183,
      data184,
      data185,
      data186,
      data187,
      data188,
      data189,
      data190,
      data191,
      data192,
      data193,
      data194,
      data195,
      data196,
      data197,
      data198,
      data199,
      data200,
      data201,
      data202,
      data203,
      data204,
      data205,
      data206,
      data207,
      data208,
      data209,
      data210,
      data211,
      data212,
      data213,
      data214,
      data215,
      data216,
      data217,
      data218,
      data219,
      data220,
      data221,
      data222,
      data223,
      data224,
      data225,
      data226,
      data227,
      data228,
      data229,
      data230,
      data231,
      data232,
      data233,
      data234,
      data235,
      data236,
      data237,
      data238,
      data239,
      data240,
      data241,
      data242,
      data243,
      data244,
      data245,
      data246,
      data247,
      data248,
      data249,
      data250,
      data251,
      data252,
      data253,
      data254,
      data255,
      data256,
      data257,
      data258,
      data259,
      data260,
      data261,
      data262,
      data263,
      data264,
      data265,
      data266,
      data267,
      data268,
      data269,
      data270,
      data271,
      data272,
      data273,
      data274,
      data275,
      data276,
      data277,
      data278,
      data279,
      data280,
      data281,
      data282,
      data283,
      data284,
      data285,
      data286,
      data287,
      data288;
  reg done_reg;
  assign done_o = (i_counter == 9 && done_reg == 0) ? 1 : 0;

  // handle with i rows and i cols

  always @(posedge clk) begin
    if (rst) begin
      i_row <= 0;
      i_col <= 0;
      done_reg <= 0;
    end else begin
      if (done_o) begin
        i_col <= (i_col == COLS - 1) ? 0 : i_col + 1;

        if (i_col == COLS - 1) begin
          if (i_row == ROWS - 1) begin
            done_reg <= 1;
          end
          i_row <= (i_row == ROWS - 1) ? 0 : i_row + 1;
        end
      end
    end
  end


  always @(posedge clk) begin
    if (rst) begin

      i_counter <= 0;
    end else begin
      if (done_i) begin
        i_counter <= (i_counter == 9) ? i_counter : i_counter + 1;
      end


    end

  end


  always @(*) begin
    if (rst) begin
      data0_o   <= 0;
      data1_o   <= 0;
      data2_o   <= 0;
      data3_o   <= 0;
      data4_o   <= 0;
      data5_o   <= 0;
      data6_o   <= 0;
      data7_o   <= 0;
      data8_o   <= 0;
      data9_o   <= 0;
      data10_o  <= 0;
      data11_o  <= 0;
      data12_o  <= 0;
      data13_o  <= 0;
      data14_o  <= 0;
      data15_o  <= 0;
      data16_o  <= 0;
      data17_o  <= 0;
      data18_o  <= 0;
      data19_o  <= 0;
      data20_o  <= 0;
      data21_o  <= 0;
      data22_o  <= 0;
      data23_o  <= 0;
      data24_o  <= 0;
      data25_o  <= 0;
      data26_o  <= 0;
      data27_o  <= 0;
      data28_o  <= 0;
      data29_o  <= 0;
      data30_o  <= 0;
      data31_o  <= 0;
      data32_o  <= 0;
      data33_o  <= 0;
      data34_o  <= 0;
      data35_o  <= 0;
      data36_o  <= 0;
      data37_o  <= 0;
      data38_o  <= 0;
      data39_o  <= 0;
      data40_o  <= 0;
      data41_o  <= 0;
      data42_o  <= 0;
      data43_o  <= 0;
      data44_o  <= 0;
      data45_o  <= 0;
      data46_o  <= 0;
      data47_o  <= 0;
      data48_o  <= 0;
      data49_o  <= 0;
      data50_o  <= 0;
      data51_o  <= 0;
      data52_o  <= 0;
      data53_o  <= 0;
      data54_o  <= 0;
      data55_o  <= 0;
      data56_o  <= 0;
      data57_o  <= 0;
      data58_o  <= 0;
      data59_o  <= 0;
      data60_o  <= 0;
      data61_o  <= 0;
      data62_o  <= 0;
      data63_o  <= 0;
      data64_o  <= 0;
      data65_o  <= 0;
      data66_o  <= 0;
      data67_o  <= 0;
      data68_o  <= 0;
      data69_o  <= 0;
      data70_o  <= 0;
      data71_o  <= 0;
      data72_o  <= 0;
      data73_o  <= 0;
      data74_o  <= 0;
      data75_o  <= 0;
      data76_o  <= 0;
      data77_o  <= 0;
      data78_o  <= 0;
      data79_o  <= 0;
      data80_o  <= 0;
      data81_o  <= 0;
      data82_o  <= 0;
      data83_o  <= 0;
      data84_o  <= 0;
      data85_o  <= 0;
      data86_o  <= 0;
      data87_o  <= 0;
      data88_o  <= 0;
      data89_o  <= 0;
      data90_o  <= 0;
      data91_o  <= 0;
      data92_o  <= 0;
      data93_o  <= 0;
      data94_o  <= 0;
      data95_o  <= 0;
      data96_o  <= 0;
      data97_o  <= 0;
      data98_o  <= 0;
      data99_o  <= 0;
      data100_o <= 0;
      data101_o <= 0;
      data102_o <= 0;
      data103_o <= 0;
      data104_o <= 0;
      data105_o <= 0;
      data106_o <= 0;
      data107_o <= 0;
      data108_o <= 0;
      data109_o <= 0;
      data110_o <= 0;
      data111_o <= 0;
      data112_o <= 0;
      data113_o <= 0;
      data114_o <= 0;
      data115_o <= 0;
      data116_o <= 0;
      data117_o <= 0;
      data118_o <= 0;
      data119_o <= 0;
      data120_o <= 0;
      data121_o <= 0;
      data122_o <= 0;
      data123_o <= 0;
      data124_o <= 0;
      data125_o <= 0;
      data126_o <= 0;
      data127_o <= 0;
      data128_o <= 0;
      data129_o <= 0;
      data130_o <= 0;
      data131_o <= 0;
      data132_o <= 0;
      data133_o <= 0;
      data134_o <= 0;
      data135_o <= 0;
      data136_o <= 0;
      data137_o <= 0;
      data138_o <= 0;
      data139_o <= 0;
      data140_o <= 0;
      data141_o <= 0;
      data142_o <= 0;
      data143_o <= 0;
      data144_o <= 0;
      data145_o <= 0;
      data146_o <= 0;
      data147_o <= 0;
      data148_o <= 0;
      data149_o <= 0;
      data150_o <= 0;
      data151_o <= 0;
      data152_o <= 0;
      data153_o <= 0;
      data154_o <= 0;
      data155_o <= 0;
      data156_o <= 0;
      data157_o <= 0;
      data158_o <= 0;
      data159_o <= 0;
      data160_o <= 0;
      data161_o <= 0;
      data162_o <= 0;
      data163_o <= 0;
      data164_o <= 0;
      data165_o <= 0;
      data166_o <= 0;
      data167_o <= 0;
      data168_o <= 0;
      data169_o <= 0;
      data170_o <= 0;
      data171_o <= 0;
      data172_o <= 0;
      data173_o <= 0;
      data174_o <= 0;
      data175_o <= 0;
      data176_o <= 0;
      data177_o <= 0;
      data178_o <= 0;
      data179_o <= 0;
      data180_o <= 0;
      data181_o <= 0;
      data182_o <= 0;
      data183_o <= 0;
      data184_o <= 0;
      data185_o <= 0;
      data186_o <= 0;
      data187_o <= 0;
      data188_o <= 0;
      data189_o <= 0;
      data190_o <= 0;
      data191_o <= 0;
      data192_o <= 0;
      data193_o <= 0;
      data194_o <= 0;
      data195_o <= 0;
      data196_o <= 0;
      data197_o <= 0;
      data198_o <= 0;
      data199_o <= 0;
      data200_o <= 0;
      data201_o <= 0;
      data202_o <= 0;
      data203_o <= 0;
      data204_o <= 0;
      data205_o <= 0;
      data206_o <= 0;
      data207_o <= 0;
      data208_o <= 0;
      data209_o <= 0;
      data210_o <= 0;
      data211_o <= 0;
      data212_o <= 0;
      data213_o <= 0;
      data214_o <= 0;
      data215_o <= 0;
      data216_o <= 0;
      data217_o <= 0;
      data218_o <= 0;
      data219_o <= 0;
      data220_o <= 0;
      data221_o <= 0;
      data222_o <= 0;
      data223_o <= 0;
      data224_o <= 0;
      data225_o <= 0;
      data226_o <= 0;
      data227_o <= 0;
      data228_o <= 0;
      data229_o <= 0;
      data230_o <= 0;
      data231_o <= 0;
      data232_o <= 0;
      data233_o <= 0;
      data234_o <= 0;
      data235_o <= 0;
      data236_o <= 0;
      data237_o <= 0;
      data238_o <= 0;
      data239_o <= 0;
      data240_o <= 0;
      data241_o <= 0;
      data242_o <= 0;
      data243_o <= 0;
      data244_o <= 0;
      data245_o <= 0;
      data246_o <= 0;
      data247_o <= 0;
      data248_o <= 0;
      data249_o <= 0;
      data250_o <= 0;
      data251_o <= 0;
      data252_o <= 0;
      data253_o <= 0;
      data254_o <= 0;
      data255_o <= 0;
      data256_o <= 0;
      data257_o <= 0;
      data258_o <= 0;
      data259_o <= 0;
      data260_o <= 0;
      data261_o <= 0;
      data262_o <= 0;
      data263_o <= 0;
      data264_o <= 0;
      data265_o <= 0;
      data266_o <= 0;
      data267_o <= 0;
      data268_o <= 0;
      data269_o <= 0;
      data270_o <= 0;
      data271_o <= 0;
      data272_o <= 0;
      data273_o <= 0;
      data274_o <= 0;
      data275_o <= 0;
      data276_o <= 0;
      data277_o <= 0;
      data278_o <= 0;
      data279_o <= 0;
      data280_o <= 0;
      data281_o <= 0;
      data282_o <= 0;
      data283_o <= 0;
      data284_o <= 0;
      data285_o <= 0;
      data286_o <= 0;
      data287_o <= 0;
      data288_o <= 0;
    end else begin
      // zero padding
      if (done_o) begin
        data0_o   <= (i_row < 9 || i_col < 9) ? 0 : data0;
        data1_o   <= (i_row < 9 || i_col < 8) ? 0 : data1;
        data2_o   <= (i_row < 9 || i_col < 7) ? 0 : data2;
        data3_o   <= (i_row < 9 || i_col < 6) ? 0 : data3;
        data4_o   <= (i_row < 9 || i_col < 5) ? 0 : data4;
        data5_o   <= (i_row < 9 || i_col < 4) ? 0 : data5;
        data6_o   <= (i_row < 9 || i_col < 3) ? 0 : data6;
        data7_o   <= (i_row < 9 || i_col < 2) ? 0 : data7;
        data8_o   <= (i_row < 9) ? 0 : data8;
        data9_o   <= (i_row < 9 || i_col > COLS - 2) ? 0 : data9;
        data10_o  <= (i_row < 9 || i_col > COLS - 3) ? 0 : data10;
        data11_o  <= (i_row < 9 || i_col > COLS - 4) ? 0 : data11;
        data12_o  <= (i_row < 9 || i_col > COLS - 5) ? 0 : data12;
        data13_o  <= (i_row < 9 || i_col > COLS - 6) ? 0 : data13;
        data14_o  <= (i_row < 9 || i_col > COLS - 7) ? 0 : data14;
        data15_o  <= (i_row < 9 || i_col > COLS - 8) ? 0 : data15;
        data16_o  <= (i_row < 9 || i_col > COLS - 9) ? 0 : data16;

        data17_o  <= (i_row < 8 || i_col < 9) ? 0 : data17;
        data18_o  <= (i_row < 8 || i_col < 8) ? 0 : data18;
        data19_o  <= (i_row < 8 || i_col < 7) ? 0 : data19;
        data20_o  <= (i_row < 8 || i_col < 6) ? 0 : data20;
        data21_o  <= (i_row < 8 || i_col < 5) ? 0 : data21;
        data22_o  <= (i_row < 8 || i_col < 4) ? 0 : data22;
        data23_o  <= (i_row < 8 || i_col < 3) ? 0 : data23;
        data24_o  <= (i_row < 8 || i_col < 2) ? 0 : data24;
        data25_o  <= (i_row < 8) ? 0 : data25;
        data26_o  <= (i_row < 8 || i_col > COLS - 2) ? 0 : data26;
        data27_o  <= (i_row < 8 || i_col > COLS - 3) ? 0 : data27;
        data28_o  <= (i_row < 8 || i_col > COLS - 4) ? 0 : data28;
        data29_o  <= (i_row < 8 || i_col > COLS - 5) ? 0 : data29;
        data30_o  <= (i_row < 8 || i_col > COLS - 6) ? 0 : data30;
        data31_o  <= (i_row < 8 || i_col > COLS - 7) ? 0 : data31;
        data32_o  <= (i_row < 8 || i_col > COLS - 8) ? 0 : data32;
        data33_o  <= (i_row < 8 || i_col > COLS - 9) ? 0 : data33;

        data34_o  <= (i_row < 7 || i_col < 9) ? 0 : data34;
        data35_o  <= (i_row < 7 || i_col < 8) ? 0 : data35;
        data36_o  <= (i_row < 7 || i_col < 7) ? 0 : data36;
        data37_o  <= (i_row < 7 || i_col < 6) ? 0 : data37;
        data38_o  <= (i_row < 7 || i_col < 5) ? 0 : data38;
        data39_o  <= (i_row < 7 || i_col < 4) ? 0 : data39;
        data40_o  <= (i_row < 7 || i_col < 3) ? 0 : data40;
        data41_o  <= (i_row < 7 || i_col < 2) ? 0 : data41;
        data42_o  <= (i_row < 7) ? 0 : data42;
        data43_o  <= (i_row < 7 || i_col > COLS - 2) ? 0 : data43;
        data44_o  <= (i_row < 7 || i_col > COLS - 3) ? 0 : data44;
        data45_o  <= (i_row < 7 || i_col > COLS - 4) ? 0 : data45;
        data46_o  <= (i_row < 7 || i_col > COLS - 5) ? 0 : data46;
        data47_o  <= (i_row < 7 || i_col > COLS - 6) ? 0 : data47;
        data48_o  <= (i_row < 7 || i_col > COLS - 7) ? 0 : data48;
        data49_o  <= (i_row < 7 || i_col > COLS - 8) ? 0 : data49;
        data50_o  <= (i_row < 7 || i_col > COLS - 9) ? 0 : data50;

        data51_o  <= (i_row < 6 || i_col < 9) ? 0 : data51;
        data52_o  <= (i_row < 6 || i_col < 8) ? 0 : data52;
        data53_o  <= (i_row < 6 || i_col < 7) ? 0 : data53;
        data54_o  <= (i_row < 6 || i_col < 6) ? 0 : data54;
        data55_o  <= (i_row < 6 || i_col < 5) ? 0 : data55;
        data56_o  <= (i_row < 6 || i_col < 4) ? 0 : data56;
        data57_o  <= (i_row < 6 || i_col < 3) ? 0 : data57;
        data58_o  <= (i_row < 6 || i_col < 2) ? 0 : data58;
        data59_o  <= (i_row < 6) ? 0 : data59;
        data60_o  <= (i_row < 6 || i_col > COLS - 2) ? 0 : data60;
        data61_o  <= (i_row < 6 || i_col > COLS - 3) ? 0 : data61;
        data62_o  <= (i_row < 6 || i_col > COLS - 4) ? 0 : data62;
        data63_o  <= (i_row < 6 || i_col > COLS - 5) ? 0 : data63;
        data64_o  <= (i_row < 6 || i_col > COLS - 6) ? 0 : data64;
        data65_o  <= (i_row < 6 || i_col > COLS - 7) ? 0 : data65;
        data66_o  <= (i_row < 6 || i_col > COLS - 8) ? 0 : data66;
        data67_o  <= (i_row < 6 || i_col > COLS - 9) ? 0 : data67;

        data68_o  <= (i_row < 5 || i_col < 9) ? 0 : data68;
        data69_o  <= (i_row < 5 || i_col < 8) ? 0 : data69;
        data70_o  <= (i_row < 5 || i_col < 7) ? 0 : data70;
        data71_o  <= (i_row < 5 || i_col < 6) ? 0 : data71;
        data72_o  <= (i_row < 5 || i_col < 5) ? 0 : data72;
        data73_o  <= (i_row < 5 || i_col < 4) ? 0 : data73;
        data74_o  <= (i_row < 5 || i_col < 3) ? 0 : data74;
        data75_o  <= (i_row < 5 || i_col < 2) ? 0 : data75;
        data76_o  <= (i_row < 5) ? 0 : data76;
        data77_o  <= (i_row < 5 || i_col > COLS - 2) ? 0 : data77;
        data78_o  <= (i_row < 5 || i_col > COLS - 3) ? 0 : data78;
        data79_o  <= (i_row < 5 || i_col > COLS - 4) ? 0 : data79;
        data80_o  <= (i_row < 5 || i_col > COLS - 5) ? 0 : data80;
        data81_o  <= (i_row < 5 || i_col > COLS - 6) ? 0 : data81;
        data82_o  <= (i_row < 5 || i_col > COLS - 7) ? 0 : data82;
        data83_o  <= (i_row < 5 || i_col > COLS - 8) ? 0 : data83;
        data84_o  <= (i_row < 5 || i_col > COLS - 9) ? 0 : data84;

        data85_o  <= (i_row < 4 || i_col < 9) ? 0 : data85;
        data86_o  <= (i_row < 4 || i_col < 8) ? 0 : data86;
        data87_o  <= (i_row < 4 || i_col < 7) ? 0 : data87;
        data88_o  <= (i_row < 4 || i_col < 6) ? 0 : data88;
        data89_o  <= (i_row < 4 || i_col < 5) ? 0 : data89;
        data90_o  <= (i_row < 4 || i_col < 4) ? 0 : data90;
        data91_o  <= (i_row < 4 || i_col < 3) ? 0 : data91;
        data92_o  <= (i_row < 4 || i_col < 2) ? 0 : data92;
        data93_o  <= (i_row < 4) ? 0 : data93;
        data94_o  <= (i_row < 4 || i_col > COLS - 2) ? 0 : data94;
        data95_o  <= (i_row < 4 || i_col > COLS - 3) ? 0 : data95;
        data96_o  <= (i_row < 4 || i_col > COLS - 4) ? 0 : data96;
        data97_o  <= (i_row < 4 || i_col > COLS - 5) ? 0 : data97;
        data98_o  <= (i_row < 4 || i_col > COLS - 6) ? 0 : data98;
        data99_o  <= (i_row < 4 || i_col > COLS - 7) ? 0 : data99;
        data100_o <= (i_row < 4 || i_col > COLS - 8) ? 0 : data100;
        data101_o <= (i_row < 4 || i_col > COLS - 9) ? 0 : data101;

        data102_o <= (i_row < 3 || i_col < 9) ? 0 : data102;
        data103_o <= (i_row < 3 || i_col < 8) ? 0 : data103;
        data104_o <= (i_row < 3 || i_col < 7) ? 0 : data104;
        data105_o <= (i_row < 3 || i_col < 6) ? 0 : data105;
        data106_o <= (i_row < 3 || i_col < 5) ? 0 : data106;
        data107_o <= (i_row < 3 || i_col < 5) ? 0 : data107;
        data108_o <= (i_row < 3 || i_col < 3) ? 0 : data108;
        data109_o <= (i_row < 3 || i_col < 2) ? 0 : data109;
        data110_o <= (i_row < 3) ? 0 : data110;
        data111_o <= (i_row < 3 || i_col > COLS - 2) ? 0 : data111;
        data112_o <= (i_row < 3 || i_col > COLS - 3) ? 0 : data112;
        data113_o <= (i_row < 3 || i_col > COLS - 4) ? 0 : data113;
        data114_o <= (i_row < 3 || i_col > COLS - 5) ? 0 : data114;
        data115_o <= (i_row < 3 || i_col > COLS - 6) ? 0 : data115;
        data116_o <= (i_row < 3 || i_col > COLS - 7) ? 0 : data116;
        data117_o <= (i_row < 3 || i_col > COLS - 8) ? 0 : data117;
        data118_o <= (i_row < 3 || i_col > COLS - 9) ? 0 : data118;

        data119_o <= (i_row < 2 || i_col < 9) ? 0 : data119;
        data120_o <= (i_row < 2 || i_col < 8) ? 0 : data120;
        data121_o <= (i_row < 2 || i_col < 7) ? 0 : data121;
        data122_o <= (i_row < 2 || i_col < 6) ? 0 : data122;
        data123_o <= (i_row < 2 || i_col < 5) ? 0 : data123;
        data124_o <= (i_row < 2 || i_col < 4) ? 0 : data124;
        data125_o <= (i_row < 2 || i_col < 3) ? 0 : data125;
        data126_o <= (i_row < 2 || i_col < 2) ? 0 : data126;
        data127_o <= (i_row < 2) ? 0 : data127;
        data128_o <= (i_row < 2 || i_col > COLS - 2) ? 0 : data128;
        data129_o <= (i_row < 2 || i_col > COLS - 3) ? 0 : data129;
        data130_o <= (i_row < 2 || i_col > COLS - 4) ? 0 : data130;
        data131_o <= (i_row < 2 || i_col > COLS - 5) ? 0 : data131;
        data132_o <= (i_row < 2 || i_col > COLS - 6) ? 0 : data132;
        data133_o <= (i_row < 2 || i_col > COLS - 7) ? 0 : data133;
        data134_o <= (i_row < 2 || i_col > COLS - 8) ? 0 : data134;
        data135_o <= (i_row < 2 || i_col > COLS - 9) ? 0 : data135;


        data136_o <= (i_col < 9) ? 0 : data136;
        data137_o <= (i_col < 8) ? 0 : data137;
        data138_o <= (i_col < 7) ? 0 : data138;
        data139_o <= (i_col < 6) ? 0 : data139;
        data140_o <= (i_col < 5) ? 0 : data140;
        data141_o <= (i_col < 4) ? 0 : data141;
        data142_o <= (i_col < 3) ? 0 : data142;
        data143_o <= (i_col < 2) ? 0 : data143;
        data144_o <= data144;
        data145_o <= (i_col > COLS - 2) ? 0 : data145;
        data146_o <= (i_col > COLS - 3) ? 0 : data146;
        data147_o <= (i_col > COLS - 4) ? 0 : data147;
        data148_o <= (i_col > COLS - 5) ? 0 : data148;
        data149_o <= (i_col > COLS - 6) ? 0 : data149;
        data150_o <= (i_col > COLS - 7) ? 0 : data150;
        data151_o <= (i_col > COLS - 8) ? 0 : data151;
        data152_o <= (i_col > COLS - 9) ? 0 : data152;


        data153_o <= (i_row > ROWS - 2 || i_col < 9) ? 0 : data153;
        data154_o <= (i_row > ROWS - 2 || i_col < 8) ? 0 : data154;
        data155_o <= (i_row > ROWS - 2 || i_col < 7) ? 0 : data155;
        data156_o <= (i_row > ROWS - 2 || i_col < 6) ? 0 : data156;
        data157_o <= (i_row > ROWS - 2 || i_col < 5) ? 0 : data157;
        data158_o <= (i_row > ROWS - 2 || i_col < 4) ? 0 : data158;
        data159_o <= (i_row > ROWS - 2 || i_col < 3) ? 0 : data159;
        data160_o <= (i_row > ROWS - 2 || i_col < 2) ? 0 : data160;
        data161_o <= (i_row > ROWS - 2) ? 0 : data161;
        data162_o <= (i_row > ROWS - 2 || i_col < COLS - 2) ? 0 : data162;
        data163_o <= (i_row > ROWS - 2 || i_col < COLS - 3) ? 0 : data163;
        data164_o <= (i_row > ROWS - 2 || i_col < COLS - 4) ? 0 : data164;
        data165_o <= (i_row > ROWS - 2 || i_col < COLS - 5) ? 0 : data165;
        data166_o <= (i_row > ROWS - 2 || i_col < COLS - 6) ? 0 : data166;
        data167_o <= (i_row > ROWS - 2 || i_col < COLS - 7) ? 0 : data167;
        data168_o <= (i_row > ROWS - 2 || i_col < COLS - 8) ? 0 : data168;
        data169_o <= (i_row > ROWS - 2 || i_col < COLS - 9) ? 0 : data169;


        data170_o <= (i_row > ROWS - 3 || i_col < 9) ? 0 : data170;
        data171_o <= (i_row > ROWS - 3 || i_col < 8) ? 0 : data171;
        data172_o <= (i_row > ROWS - 3 || i_col < 7) ? 0 : data172;
        data173_o <= (i_row > ROWS - 3 || i_col < 6) ? 0 : data173;
        data174_o <= (i_row > ROWS - 3 || i_col < 5) ? 0 : data174;
        data175_o <= (i_row > ROWS - 3 || i_col < 4) ? 0 : data175;
        data176_o <= (i_row > ROWS - 3 || i_col < 3) ? 0 : data176;
        data177_o <= (i_row > ROWS - 3 || i_col < 2) ? 0 : data177;
        data178_o <= (i_row > ROWS - 3) ? 0 : data178;
        data179_o <= (i_row > ROWS - 3 || i_col < COLS - 2) ? 0 : data179;
        data180_o <= (i_row > ROWS - 3 || i_col < COLS - 3) ? 0 : data180;
        data181_o <= (i_row > ROWS - 3 || i_col < COLS - 4) ? 0 : data181;
        data182_o <= (i_row > ROWS - 3 || i_col < COLS - 5) ? 0 : data182;
        data183_o <= (i_row > ROWS - 3 || i_col < COLS - 6) ? 0 : data183;
        data184_o <= (i_row > ROWS - 3 || i_col < COLS - 7) ? 0 : data184;
        data185_o <= (i_row > ROWS - 3 || i_col < COLS - 8) ? 0 : data185;
        data186_o <= (i_row > ROWS - 3 || i_col < COLS - 9) ? 0 : data186;

        data187_o <= (i_row > ROWS - 4 || i_col < 9) ? 0 : data187;
        data188_o <= (i_row > ROWS - 4 || i_col < 8) ? 0 : data188;
        data189_o <= (i_row > ROWS - 4 || i_col < 7) ? 0 : data189;
        data190_o <= (i_row > ROWS - 4 || i_col < 6) ? 0 : data190;
        data191_o <= (i_row > ROWS - 4 || i_col < 5) ? 0 : data191;
        data192_o <= (i_row > ROWS - 4 || i_col < 4) ? 0 : data192;
        data193_o <= (i_row > ROWS - 4 || i_col < 3) ? 0 : data193;
        data194_o <= (i_row > ROWS - 4 || i_col < 2) ? 0 : data194;
        data195_o <= (i_row > ROWS - 4) ? 0 : data195;
        data196_o <= (i_row > ROWS - 4 || i_col < COLS - 2) ? 0 : data196;
        data197_o <= (i_row > ROWS - 4 || i_col < COLS - 3) ? 0 : data197;
        data198_o <= (i_row > ROWS - 4 || i_col < COLS - 4) ? 0 : data198;
        data199_o <= (i_row > ROWS - 4 || i_col < COLS - 5) ? 0 : data199;
        data200_o <= (i_row > ROWS - 4 || i_col < COLS - 6) ? 0 : data200;
        data201_o <= (i_row > ROWS - 4 || i_col < COLS - 7) ? 0 : data201;
        data202_o <= (i_row > ROWS - 4 || i_col < COLS - 8) ? 0 : data202;
        data203_o <= (i_row > ROWS - 4 || i_col < COLS - 9) ? 0 : data203;


        data204_o <= (i_row > ROWS - 5 || i_col < 9) ? 0 : data204;
        data205_o <= (i_row > ROWS - 5 || i_col < 8) ? 0 : data205;
        data206_o <= (i_row > ROWS - 5 || i_col < 7) ? 0 : data206;
        data207_o <= (i_row > ROWS - 5 || i_col < 6) ? 0 : data207;
        data208_o <= (i_row > ROWS - 5 || i_col < 5) ? 0 : data208;
        data209_o <= (i_row > ROWS - 5 || i_col < 4) ? 0 : data209;
        data210_o <= (i_row > ROWS - 5 || i_col < 3) ? 0 : data210;
        data211_o <= (i_row > ROWS - 5 || i_col < 2) ? 0 : data211;
        data212_o <= (i_row > ROWS - 5) ? 0 : data212;
        data213_o <= (i_row > ROWS - 5 || i_col < COLS - 2) ? 0 : data213;
        data214_o <= (i_row > ROWS - 5 || i_col < COLS - 3) ? 0 : data214;
        data215_o <= (i_row > ROWS - 5 || i_col < COLS - 4) ? 0 : data215;
        data216_o <= (i_row > ROWS - 5 || i_col < COLS - 5) ? 0 : data216;
        data217_o <= (i_row > ROWS - 5 || i_col < COLS - 6) ? 0 : data217;
        data218_o <= (i_row > ROWS - 5 || i_col < COLS - 7) ? 0 : data218;
        data219_o <= (i_row > ROWS - 5 || i_col < COLS - 8) ? 0 : data219;
        data220_o <= (i_row > ROWS - 5 || i_col < COLS - 9) ? 0 : data220;

        data221_o <= (i_row > ROWS - 6 || i_col < 9) ? 0 : data221;
        data222_o <= (i_row > ROWS - 6 || i_col < 8) ? 0 : data222;
        data223_o <= (i_row > ROWS - 6 || i_col < 7) ? 0 : data223;
        data224_o <= (i_row > ROWS - 6 || i_col < 6) ? 0 : data224;
        data225_o <= (i_row > ROWS - 6 || i_col < 5) ? 0 : data225;
        data226_o <= (i_row > ROWS - 6 || i_col < 4) ? 0 : data226;
        data227_o <= (i_row > ROWS - 6 || i_col < 3) ? 0 : data227;
        data228_o <= (i_row > ROWS - 6 || i_col < 2) ? 0 : data228;
        data229_o <= (i_row > ROWS - 6) ? 0 : data229;
        data230_o <= (i_row > ROWS - 6 || i_col < COLS - 2) ? 0 : data230;
        data231_o <= (i_row > ROWS - 6 || i_col < COLS - 3) ? 0 : data231;
        data232_o <= (i_row > ROWS - 6 || i_col < COLS - 4) ? 0 : data232;
        data233_o <= (i_row > ROWS - 6 || i_col < COLS - 5) ? 0 : data233;
        data234_o <= (i_row > ROWS - 6 || i_col < COLS - 6) ? 0 : data234;
        data235_o <= (i_row > ROWS - 6 || i_col < COLS - 7) ? 0 : data235;
        data236_o <= (i_row > ROWS - 6 || i_col < COLS - 8) ? 0 : data236;
        data237_o <= (i_row > ROWS - 6 || i_col < COLS - 9) ? 0 : data237;

        data238_o <= (i_row > ROWS - 7 || i_col < 9) ? 0 : data238;
        data239_o <= (i_row > ROWS - 7 || i_col < 8) ? 0 : data239;
        data240_o <= (i_row > ROWS - 7 || i_col < 7) ? 0 : data240;
        data241_o <= (i_row > ROWS - 7 || i_col < 6) ? 0 : data241;
        data242_o <= (i_row > ROWS - 7 || i_col < 5) ? 0 : data242;
        data243_o <= (i_row > ROWS - 7 || i_col < 4) ? 0 : data243;
        data244_o <= (i_row > ROWS - 7 || i_col < 3) ? 0 : data244;
        data245_o <= (i_row > ROWS - 7 || i_col < 2) ? 0 : data245;
        data246_o <= (i_row > ROWS - 7) ? 0 : data246;
        data247_o <= (i_row > ROWS - 7 || i_col < COLS - 2) ? 0 : data247;
        data248_o <= (i_row > ROWS - 7 || i_col < COLS - 3) ? 0 : data248;
        data249_o <= (i_row > ROWS - 7 || i_col < COLS - 4) ? 0 : data249;
        data250_o <= (i_row > ROWS - 7 || i_col < COLS - 5) ? 0 : data250;
        data251_o <= (i_row > ROWS - 7 || i_col < COLS - 6) ? 0 : data251;
        data252_o <= (i_row > ROWS - 7 || i_col < COLS - 7) ? 0 : data252;
        data253_o <= (i_row > ROWS - 7 || i_col < COLS - 8) ? 0 : data253;
        data254_o <= (i_row > ROWS - 7 || i_col < COLS - 9) ? 0 : data254;

        data255_o <= (i_row > ROWS - 8 || i_col < 9) ? 0 : data255;
        data256_o <= (i_row > ROWS - 8 || i_col < 8) ? 0 : data256;
        data257_o <= (i_row > ROWS - 8 || i_col < 7) ? 0 : data257;
        data258_o <= (i_row > ROWS - 8 || i_col < 6) ? 0 : data258;
        data259_o <= (i_row > ROWS - 8 || i_col < 5) ? 0 : data259;
        data260_o <= (i_row > ROWS - 8 || i_col < 4) ? 0 : data260;
        data261_o <= (i_row > ROWS - 8 || i_col < 3) ? 0 : data261;
        data262_o <= (i_row > ROWS - 8 || i_col < 2) ? 0 : data262;
        data263_o <= (i_row > ROWS - 8) ? 0 : data263;
        data264_o <= (i_row > ROWS - 8 || i_col < COLS - 2) ? 0 : data264;
        data265_o <= (i_row > ROWS - 8 || i_col < COLS - 3) ? 0 : data265;
        data266_o <= (i_row > ROWS - 8 || i_col < COLS - 4) ? 0 : data266;
        data267_o <= (i_row > ROWS - 8 || i_col < COLS - 5) ? 0 : data267;
        data268_o <= (i_row > ROWS - 8 || i_col < COLS - 6) ? 0 : data268;
        data269_o <= (i_row > ROWS - 8 || i_col < COLS - 7) ? 0 : data269;
        data270_o <= (i_row > ROWS - 8 || i_col < COLS - 8) ? 0 : data270;
        data271_o <= (i_row > ROWS - 8 || i_col < COLS - 9) ? 0 : data271;

        data272_o <= (i_row > ROWS - 9 || i_col < 9) ? 0 : data272;
        data273_o <= (i_row > ROWS - 9 || i_col < 8) ? 0 : data273;
        data274_o <= (i_row > ROWS - 9 || i_col < 7) ? 0 : data274;
        data275_o <= (i_row > ROWS - 9 || i_col < 6) ? 0 : data275;
        data276_o <= (i_row > ROWS - 9 || i_col < 5) ? 0 : data276;
        data277_o <= (i_row > ROWS - 9 || i_col < 4) ? 0 : data277;
        data278_o <= (i_row > ROWS - 9 || i_col < 3) ? 0 : data278;
        data279_o <= (i_row > ROWS - 9 || i_col < 2) ? 0 : data279;
        data280_o <= (i_row > ROWS - 9) ? 0 : data280;
        data281_o <= (i_row > ROWS - 9 || i_col < COLS - 2) ? 0 : data281;
        data282_o <= (i_row > ROWS - 9 || i_col < COLS - 3) ? 0 : data282;
        data283_o <= (i_row > ROWS - 9 || i_col < COLS - 4) ? 0 : data283;
        data284_o <= (i_row > ROWS - 9 || i_col < COLS - 5) ? 0 : data284;
        data285_o <= (i_row > ROWS - 9 || i_col < COLS - 6) ? 0 : data285;
        data286_o <= (i_row > ROWS - 9 || i_col < COLS - 7) ? 0 : data286;
        data287_o <= (i_row > ROWS - 9 || i_col < COLS - 8) ? 0 : data287;
        data288_o <= (i_row > ROWS - 9 || i_col < COLS - 9) ? 0 : data288;

      end
    end
  end

  always @(posedge clk) begin
    if (rst) begin
      data0   <= 0;
      data1   <= 0;
      data2   <= 0;
      data3   <= 0;
      data4   <= 0;
      data5   <= 0;
      data6   <= 0;
      data7   <= 0;
      data8   <= 0;
      data9   <= 0;
      data10  <= 0;
      data11  <= 0;
      data12  <= 0;
      data13  <= 0;
      data14  <= 0;
      data15  <= 0;
      data16  <= 0;
      data17  <= 0;
      data18  <= 0;
      data19  <= 0;
      data20  <= 0;
      data21  <= 0;
      data22  <= 0;
      data23  <= 0;
      data24  <= 0;
      data25  <= 0;
      data26  <= 0;
      data27  <= 0;
      data28  <= 0;
      data29  <= 0;
      data30  <= 0;
      data31  <= 0;
      data32  <= 0;
      data33  <= 0;
      data34  <= 0;
      data35  <= 0;
      data36  <= 0;
      data37  <= 0;
      data38  <= 0;
      data39  <= 0;
      data40  <= 0;
      data41  <= 0;
      data42  <= 0;
      data43  <= 0;
      data44  <= 0;
      data45  <= 0;
      data46  <= 0;
      data47  <= 0;
      data48  <= 0;
      data49  <= 0;
      data50  <= 0;
      data51  <= 0;
      data52  <= 0;
      data53  <= 0;
      data54  <= 0;
      data55  <= 0;
      data56  <= 0;
      data57  <= 0;
      data58  <= 0;
      data59  <= 0;
      data60  <= 0;
      data61  <= 0;
      data62  <= 0;
      data63  <= 0;
      data64  <= 0;
      data65  <= 0;
      data66  <= 0;
      data67  <= 0;
      data68  <= 0;
      data69  <= 0;
      data70  <= 0;
      data71  <= 0;
      data72  <= 0;
      data73  <= 0;
      data74  <= 0;
      data75  <= 0;
      data76  <= 0;
      data77  <= 0;
      data78  <= 0;
      data79  <= 0;
      data80  <= 0;
      data81  <= 0;
      data82  <= 0;
      data83  <= 0;
      data84  <= 0;
      data85  <= 0;
      data86  <= 0;
      data87  <= 0;
      data88  <= 0;
      data89  <= 0;
      data90  <= 0;
      data91  <= 0;
      data92  <= 0;
      data93  <= 0;
      data94  <= 0;
      data95  <= 0;
      data96  <= 0;
      data97  <= 0;
      data98  <= 0;
      data99  <= 0;
      data100 <= 0;
      data101 <= 0;
      data102 <= 0;
      data103 <= 0;
      data104 <= 0;
      data105 <= 0;
      data106 <= 0;
      data107 <= 0;
      data108 <= 0;
      data109 <= 0;
      data110 <= 0;
      data111 <= 0;
      data112 <= 0;
      data113 <= 0;
      data114 <= 0;
      data115 <= 0;
      data116 <= 0;
      data117 <= 0;
      data118 <= 0;
      data119 <= 0;
      data120 <= 0;
      data121 <= 0;
      data122 <= 0;
      data123 <= 0;
      data124 <= 0;
      data125 <= 0;
      data126 <= 0;
      data127 <= 0;
      data128 <= 0;
      data129 <= 0;
      data130 <= 0;
      data131 <= 0;
      data132 <= 0;
      data133 <= 0;
      data134 <= 0;
      data135 <= 0;
      data136 <= 0;
      data137 <= 0;
      data138 <= 0;
      data139 <= 0;
      data140 <= 0;
      data141 <= 0;
      data142 <= 0;
      data143 <= 0;
      data144 <= 0;
      data145 <= 0;
      data146 <= 0;
      data147 <= 0;
      data148 <= 0;
      data149 <= 0;
      data150 <= 0;
      data151 <= 0;
      data152 <= 0;
      data153 <= 0;
      data154 <= 0;
      data155 <= 0;
      data156 <= 0;
      data157 <= 0;
      data158 <= 0;
      data159 <= 0;
      data160 <= 0;
      data161 <= 0;
      data162 <= 0;
      data163 <= 0;
      data164 <= 0;
      data165 <= 0;
      data166 <= 0;
      data167 <= 0;
      data168 <= 0;
      data169 <= 0;
      data170 <= 0;
      data171 <= 0;
      data172 <= 0;
      data173 <= 0;
      data174 <= 0;
      data175 <= 0;
      data176 <= 0;
      data177 <= 0;
      data178 <= 0;
      data179 <= 0;
      data180 <= 0;
      data181 <= 0;
      data182 <= 0;
      data183 <= 0;
      data184 <= 0;
      data185 <= 0;
      data186 <= 0;
      data187 <= 0;
      data188 <= 0;
      data189 <= 0;
      data190 <= 0;
      data191 <= 0;
      data192 <= 0;
      data193 <= 0;
      data194 <= 0;
      data195 <= 0;
      data196 <= 0;
      data197 <= 0;
      data198 <= 0;
      data199 <= 0;
      data200 <= 0;
      data201 <= 0;
      data202 <= 0;
      data203 <= 0;
      data204 <= 0;
      data205 <= 0;
      data206 <= 0;
      data207 <= 0;
      data208 <= 0;
      data209 <= 0;
      data210 <= 0;
      data211 <= 0;
      data212 <= 0;
      data213 <= 0;
      data214 <= 0;
      data215 <= 0;
      data216 <= 0;
      data217 <= 0;
      data218 <= 0;
      data219 <= 0;
      data220 <= 0;
      data221 <= 0;
      data222 <= 0;
      data223 <= 0;
      data224 <= 0;
      data225 <= 0;
      data226 <= 0;
      data227 <= 0;
      data228 <= 0;
      data229 <= 0;
      data230 <= 0;
      data231 <= 0;
      data232 <= 0;
      data233 <= 0;
      data234 <= 0;
      data235 <= 0;
      data236 <= 0;
      data237 <= 0;
      data238 <= 0;
      data239 <= 0;
      data240 <= 0;
      data241 <= 0;
      data242 <= 0;
      data243 <= 0;
      data244 <= 0;
      data245 <= 0;
      data246 <= 0;
      data247 <= 0;
      data248 <= 0;
      data249 <= 0;
      data250 <= 0;
      data251 <= 0;
      data252 <= 0;
      data253 <= 0;
      data254 <= 0;
      data255 <= 0;
      data256 <= 0;
      data257 <= 0;
      data258 <= 0;
      data259 <= 0;
      data260 <= 0;
      data261 <= 0;
      data262 <= 0;
      data263 <= 0;
      data264 <= 0;
      data265 <= 0;
      data266 <= 0;
      data267 <= 0;
      data268 <= 0;
      data269 <= 0;
      data270 <= 0;
      data271 <= 0;
      data272 <= 0;
      data273 <= 0;
      data274 <= 0;
      data275 <= 0;
      data276 <= 0;
      data277 <= 0;
      data278 <= 0;
      data279 <= 0;
      data280 <= 0;
      data281 <= 0;
      data282 <= 0;
      data283 <= 0;
      data284 <= 0;
      data285 <= 0;
      data286 <= 0;
      data287 <= 0;
      data288 <= 0;
    end else begin
      // d7 d6 d5 d4 d3 d2 d1
      if (done_i) begin
        data0   <= data1;
        data1   <= data2;
        data2   <= data3;
        data3   <= data4;
        data4   <= data5;
        data5   <= data6;
        data6   <= data7;
        data7   <= data8;
        data8   <= data9;
        data9   <= data10;
        data10  <= data11;
        data11  <= data12;
        data12  <= data13;
        data13  <= data14;
        data14  <= data15;
        data15  <= data16;
        data16  <= data16_i;

        data17  <= data18;
        data18  <= data19;
        data19  <= data20;
        data20  <= data21;
        data21  <= data22;
        data22  <= data23;
        data23  <= data24;
        data24  <= data25;
        data25  <= data26;
        data26  <= data27;
        data27  <= data28;
        data28  <= data29;
        data29  <= data30;
        data30  <= data31;
        data31  <= data32;
        data32  <= data33;
        data33  <= data15_i;


        data51  <= data52;
        data52  <= data53;
        data53  <= data54;
        data54  <= data55;
        data55  <= data56;
        data56  <= data57;
        data57  <= data58;
        data58  <= data59;
        data59  <= data60;
        data60  <= data61;
        data61  <= data62;
        data62  <= data63;
        data63  <= data64;
        data64  <= data65;
        data65  <= data66;
        data66  <= data67;
        data67  <= data14_i;


        data51  <= data52;
        data52  <= data53;
        data53  <= data54;
        data54  <= data55;
        data55  <= data56;
        data56  <= data57;
        data57  <= data58;
        data58  <= data59;
        data59  <= data60;
        data60  <= data61;
        data61  <= data62;
        data62  <= data63;
        data63  <= data64;
        data64  <= data65;
        data65  <= data66;
        data66  <= data67;
        data67  <= data13_i;


        data68  <= data69;
        data69  <= data70;
        data70  <= data71;
        data71  <= data72;
        data72  <= data73;
        data73  <= data74;
        data74  <= data75;
        data75  <= data76;
        data76  <= data77;
        data77  <= data78;
        data78  <= data79;
        data79  <= data80;
        data80  <= data81;
        data81  <= data82;
        data82  <= data83;
        data83  <= data84;
        data84  <= data12_i;

        data85  <= data86;
        data86  <= data87;
        data87  <= data88;
        data88  <= data89;
        data89  <= data90;
        data90  <= data91;
        data91  <= data92;
        data92  <= data93;
        data93  <= data94;
        data94  <= data95;
        data95  <= data96;
        data96  <= data97;
        data97  <= data98;
        data98  <= data99;
        data99  <= data100;
        data100 <= data101;
        data101 <= data11_i;

        data102 <= data103;
        data103 <= data104;
        data104 <= data105;
        data105 <= data106;
        data106 <= data107;
        data107 <= data108;
        data108 <= data109;
        data109 <= data110;
        data110 <= data111;
        data111 <= data112;
        data112 <= data113;
        data113 <= data114;
        data114 <= data115;
        data115 <= data116;
        data116 <= data117;
        data117 <= data118;
        data118 <= data10_i;

        data119 <= data120;
        data120 <= data121;
        data121 <= data122;
        data122 <= data123;
        data123 <= data124;
        data124 <= data125;
        data125 <= data126;
        data126 <= data127;
        data127 <= data128;
        data128 <= data129;
        data129 <= data130;
        data130 <= data131;
        data131 <= data132;
        data132 <= data133;
        data133 <= data134;
        data134 <= data135;
        data135 <= data9_i;

        data136 <= data137;
        data137 <= data138;
        data138 <= data139;
        data139 <= data140;
        data140 <= data141;
        data141 <= data142;
        data142 <= data143;
        data143 <= data144;
        data144 <= data145;
        data145 <= data146;
        data146 <= data147;
        data147 <= data148;
        data148 <= data149;
        data149 <= data150;
        data150 <= data151;
        data151 <= data152;
        data152 <= data8_i;

        data153 <= data154;
        data154 <= data155;
        data155 <= data156;
        data156 <= data157;
        data157 <= data158;
        data158 <= data159;
        data159 <= data160;
        data160 <= data161;
        data161 <= data162;
        data162 <= data163;
        data163 <= data164;
        data164 <= data165;
        data165 <= data166;
        data166 <= data167;
        data167 <= data168;
        data168 <= data169;
        data169 <= data7_i;

        data170 <= data171;
        data171 <= data172;
        data172 <= data173;
        data173 <= data174;
        data174 <= data175;
        data175 <= data176;
        data176 <= data177;
        data177 <= data178;
        data178 <= data179;
        data179 <= data180;
        data180 <= data181;
        data181 <= data182;
        data182 <= data183;
        data183 <= data184;
        data184 <= data185;
        data185 <= data186;
        data186 <= data6_i;

        data187 <= data188;
        data188 <= data189;
        data189 <= data190;
        data190 <= data191;
        data191 <= data192;
        data192 <= data193;
        data193 <= data194;
        data194 <= data195;
        data195 <= data196;
        data196 <= data197;
        data197 <= data198;
        data198 <= data199;
        data199 <= data200;
        data200 <= data201;
        data201 <= data202;
        data202 <= data203;
        data203 <= data5_i;

        data204 <= data205;
        data205 <= data206;
        data206 <= data207;
        data207 <= data208;
        data208 <= data209;
        data209 <= data210;
        data210 <= data211;
        data211 <= data212;
        data212 <= data213;
        data213 <= data214;
        data214 <= data215;
        data215 <= data216;
        data216 <= data217;
        data217 <= data218;
        data218 <= data219;
        data219 <= data220;
        data220 <= data4_i;

        data221 <= data222;
        data222 <= data223;
        data223 <= data224;
        data224 <= data225;
        data225 <= data226;
        data226 <= data227;
        data227 <= data228;
        data228 <= data229;
        data229 <= data230;
        data230 <= data231;
        data231 <= data232;
        data232 <= data233;
        data233 <= data234;
        data234 <= data235;
        data235 <= data236;
        data236 <= data237;
        data237 <= data3_i;

        data238 <= data239;
        data239 <= data240;
        data240 <= data241;
        data241 <= data242;
        data242 <= data243;
        data243 <= data244;
        data244 <= data245;
        data245 <= data246;
        data246 <= data247;
        data247 <= data248;
        data248 <= data249;
        data249 <= data250;
        data250 <= data251;
        data251 <= data252;
        data252 <= data253;
        data253 <= data254;
        data254 <= data2_i;

        data255 <= data256;
        data256 <= data257;
        data257 <= data258;
        data258 <= data259;
        data259 <= data260;
        data260 <= data261;
        data261 <= data262;
        data262 <= data263;
        data263 <= data264;
        data264 <= data265;
        data265 <= data266;
        data266 <= data267;
        data267 <= data268;
        data268 <= data269;
        data269 <= data270;
        data270 <= data271;
        data271 <= data1_i;

        data272 <= data273;
        data273 <= data274;
        data274 <= data275;
        data275 <= data276;
        data276 <= data277;
        data277 <= data278;
        data278 <= data279;
        data279 <= data280;
        data280 <= data281;
        data281 <= data282;
        data282 <= data283;
        data283 <= data284;
        data284 <= data285;
        data285 <= data286;
        data286 <= data287;
        data287 <= data288;
        data288 <= data0_i;

      end

    end
  end

endmodule
