module Window_buffer_9x9 #(parameter COLS = 11,
                           parameter ROWS = 11)
                          (input clk,
                           input rst_n,
                           input done_i,
                           input[7:0] S1_i,
                           S2_i,
                           S3_i,
                           S4_i,
                           S5_i,
                           S6_i,
                           S7_i,
                           S8_i,
                           S9_i,
                           output[7:0] S1_o,
                           S2_o,
                           S3_o,
                           S4_o,
                           S5_o,
                           S6_o,
                           S7_o,
                           S8_o,
                           S9_o,
                           S10_o,
                           S11_o,
                           S12_o,
                           S13_o,
                           S14_o,
                           S15_o,
                           S16_o,
                           S17_o,
                           S18_o,
                           S19_o,
                           S20_o,
                           S21_o,
                           S22_o,
                           S23_o,
                           S24_o,
                           S25_o,
                           S26_o,
                           S27_o,
                           S28_o,
                           S29_o,
                           S30_o,
                           S31_o,
                           S32_o,
                           S33_o,
                           S34_o,
                           S35_o,
                           S36_o,
                           S37_o,
                           S38_o,
                           S39_o,
                           S40_o,
                           S41_o,
                           S42_o,
                           S43_o,
                           S44_o,
                           S45_o,
                           S46_o,
                           S47_o,
                           S48_o,
                           S49_o,
                           S50_o,
                           S51_o,
                           S52_o,
                           S53_o,
                           S54_o,
                           S55_o,
                           S56_o,
                           S57_o,
                           S58_o,
                           S59_o,
                           S60_o,
                           S61_o,
                           S62_o,
                           S63_o,
                           S64_o,
                           S65_o,
                           S66_o,
                           S67_o,
                           S68_o,
                           S69_o,
                           S70_o,
                           S71_o,
                           S72_o,
                           S73_o,
                           S74_o,
                           S75_o,
                           S76_o,
                           S77_o,
                           S78_o,
                           S79_o,
                           S80_o,
                           S81_o,
                           output done_o,
                           output progress_done_o);
    wire i_row_eq_max, i_col_eq_max, i_col_ge_threshold;
    wire count_en;
    Window_buffer_9x9_controller WINDOW_BUFFER_9X9_CONTROLLER(
    .clk(clk),
    .rst_n(rst_n),
    .done_i(done_i),
    .i_row_eq_max(i_row_eq_max),
    .i_col_eq_max(i_col_eq_max),
    .i_col_ge_threshold(i_col_ge_threshold),
    .count_en(count_en),
    .progress_done(progress_done_o),
    .done_o(done_o));
    
    Window_buffer_9x9_datapath #(.COLS(COLS),
    .ROWS(ROWS))
    WINDOW_BUFFER_9X9_DATAPATH
    (
    .clk(clk),
    .rst_n(rst_n),
    .count_en(count_en),
    .S1_i(S1_i),
    .S2_i(S2_i),
    .S3_i(S3_i),
    .S4_i(S4_i),
    .S5_i(S5_i),
    .S6_i(S6_i),
    .S7_i(S7_i),
    .S8_i(S8_i),
    .S9_i(S9_i),
    .i_row_eq_max(i_row_eq_max),
    .S1_o(S1_o),
    .S2_o(S2_o),
    .S3_o(S3_o),
    .S4_o(S4_o),
    .S5_o(S5_o),
    .S6_o(S6_o),
    .S7_o(S7_o),
    .S8_o(S8_o),
    .S9_o(S9_o),
    .S10_o(S10_o),
    .S11_o(S11_o),
    .S12_o(S12_o),
    .S13_o(S13_o),
    .S14_o(S14_o),
    .S15_o(S15_o),
    .S16_o(S16_o),
    .S17_o(S17_o),
    .S18_o(S18_o),
    .S19_o(S19_o),
    .S20_o(S20_o),
    .S21_o(S21_o),
    .S22_o(S22_o),
    .S23_o(S23_o),
    .S24_o(S24_o),
    .S25_o(S25_o),
    .S26_o(S26_o),
    .S27_o(S27_o),
    .S28_o(S28_o),
    .S29_o(S29_o),
    .S30_o(S30_o),
    .S31_o(S31_o),
    .S32_o(S32_o),
    .S33_o(S33_o),
    .S34_o(S34_o),
    .S35_o(S35_o),
    .S36_o(S36_o),
    .S37_o(S37_o),
    .S38_o(S38_o),
    .S39_o(S39_o),
    .S40_o(S40_o),
    .S41_o(S41_o),
    .S42_o(S42_o),
    .S43_o(S43_o),
    .S44_o(S44_o),
    .S45_o(S45_o),
    .S46_o(S46_o),
    .S47_o(S47_o),
    .S48_o(S48_o),
    .S49_o(S49_o),
    .S50_o(S50_o),
    .S51_o(S51_o),
    .S52_o(S52_o),
    .S53_o(S53_o),
    .S54_o(S54_o),
    .S55_o(S55_o),
    .S56_o(S56_o),
    .S57_o(S57_o),
    .S58_o(S58_o),
    .S59_o(S59_o),
    .S60_o(S60_o),
    .S61_o(S61_o),
    .S62_o(S62_o),
    .S63_o(S63_o),
    .S64_o(S64_o),
    .S65_o(S65_o),
    .S66_o(S66_o),
    .S67_o(S67_o),
    .S68_o(S68_o),
    .S69_o(S69_o),
    .S70_o(S70_o),
    .S71_o(S71_o),
    .S72_o(S72_o),
    .S73_o(S73_o),
    .S74_o(S74_o),
    .S75_o(S75_o),
    .S76_o(S76_o),
    .S77_o(S77_o),
    .S78_o(S78_o),
    .S79_o(S79_o),
    .S80_o(S80_o),
    .S81_o(S81_o),
    .i_col_eq_max(i_col_eq_max),
    .i_col_ge_threshold(i_col_ge_threshold));
    
endmodule
