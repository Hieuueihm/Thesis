module Window_buffer_3x3_controller(input clk,
                                    input rst,
                                    input done_i,
                                    input [9:0] i_counter,
                                    input i_row_eq_max,
                                    output count_en,
                                    );
    
    
endmodule
