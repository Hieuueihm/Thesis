module Median_filter_5x5 #(parameter ROWS = 7,
                           parameter COLS = 7)
                          (input clk,
                           input rst_n,
                           input done_i,
                           input [7:0] d0_i,
                           input [7:0] d1_i,
                           input [7:0] d2_i,
                           input [7:0] d3_i,
                           input [7:0] d4_i,
                           output [7:0] median_o,
                           output done_o);
    wire [7:0]
    data0,
    data1,
    data2,
    data3,
    data4,
    data5,
    data6,
    data7,
    data8,
    data9,
    data10,
    data11,
    data12,
    data13,
    data14,
    data15,
    data16,
    data17,
    data18,
    data19,
    data20,
    data21,
    data22,
    data23,
    data24;
    wire done_o_modulate;
    Data_modulate_5x5 #(
    .ROWS(ROWS),
    .COLS(COLS)
    ) MEDIAN_5x5_DATA_MODULATE (
    .clk(clk),
    .rst_n(rst_n),
    .d0_i(d0_i),  // 99
    .d1_i(d1_i),  // 8
    .d2_i(d2_i),  // 7
    .d3_i(d3_i),
    .d4_i(d4_i),
    // d5 d4 d3
    .done_i(done_i),
    .d0_o(data0),
    .d1_o(data1),
    .d2_o(data2),
    .d3_o(data3),
    .d4_o(data4),
    .d5_o(data5),
    .d6_o(data6),
    .d7_o(data7),
    .d8_o(data8),
    .d9_o(data9),
    .d10_o(data10),
    .d11_o(data11),
    .d12_o(data12),
    .d13_o(data13),
    .d14_o(data14),
    .d15_o(data15),
    .d16_o(data16),
    .d17_o(data17),
    .d18_o(data18),
    .d19_o(data19),
    .d20_o(data20),
    .d21_o(data21),
    .d22_o(data22),
    .d23_o(data23),
    .d24_o(data24),
    .done_o(done_o_modulate)
    
    );
    
    Median_filter_5x5_calc MEDIAN_5X5_CALC (
    .clk(clk),
    .rst_n(rst_n),
    .done_i(done_o_modulate),
    .S1(data0),
    .S2(data1),
    .S3(data2),
    .S4(data3),
    .S5(data4),
    .S6(data5),
    .S7(data6),
    .S8(data7),
    .S9(data8),
    .S10(data9),
    .S11(data10),
    .S12(data11),
    .S13(data12),
    .S14(data13),
    .S15(data14),
    .S16(data15),
    .S17(data16),
    .S18(data17),
    .S19(data18),
    .S20(data19),
    .S21(data20),
    .S22(data21),
    .S23(data22),
    .S24(data23),
    .S25(data24),
    .median_o(median_o),
    .done_o(done_o)
    );
    
    
    
endmodule
