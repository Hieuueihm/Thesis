module data_modulate_7x7 #(
    parameter ROWS = 7,
    parameter COLS = 7
) (
    input clk,
    input rst_n,
    input [7:0] d0_i,
    input [7:0] d1_i,
    input [7:0] d2_i,
    input [7:0] d3_i,
    input [7:0] d4_i,
    input [7:0] d5_i,
    input [7:0] d6_i,
    input done_i,
    output [7:0] d0_o,
    output [7:0] d1_o,
    output [7:0] d2_o,
    output [7:0] d3_o,
    output [7:0] d4_o,
    output [7:0] d5_o,
    output [7:0] d6_o,
    output [7:0] d7_o,
    output [7:0] d8_o,
    output [7:0] d9_o,
    output [7:0] d10_o,
    output [7:0] d11_o,
    output [7:0] d12_o,
    output [7:0] d13_o,
    output [7:0] d14_o,
    output [7:0] d15_o,
    output [7:0] d16_o,
    output [7:0] d17_o,
    output [7:0] d18_o,
    output [7:0] d19_o,
    output [7:0] d20_o,
    output [7:0] d21_o,
    output [7:0] d22_o,
    output [7:0] d23_o,
    output [7:0] d24_o,
    output [7:0] d25_o,
    output [7:0] d26_o,
    output [7:0] d27_o,
    output [7:0] d28_o,
    output [7:0] d29_o,
    output [7:0] d30_o,
    output [7:0] d31_o,
    output [7:0] d32_o,
    output [7:0] d33_o,
    output [7:0] d34_o,
    output [7:0] d35_o,
    output [7:0] d36_o,
    output [7:0] d37_o,
    output [7:0] d38_o,
    output [7:0] d39_o,
    output [7:0] d40_o,
    output [7:0] d41_o,
    output [7:0] d42_o,
    output [7:0] d43_o,
    output [7:0] d44_o,
    output [7:0] d45_o,
    output [7:0] d46_o,
    output [7:0] d47_o,
    output [7:0] d48_o,
    output done_o
);

  wire finish_en;
  wire o_en;
  wire count_en;
  wire reset_en;
  wire padding_fi;
  data_modulate_7x7_controller CONTROLLER_7x7 (
      .rst_n(rst_n),
      .clk(clk),
      .done_i(done_i),
      .padding_fi(padding_fi),
      .finish_en(finish_en),
      .o_en(o_en),
      .o_valid(done_o),
      .count_en(count_en),
      .reset_en(reset_en)
  );
  data_modulate_7x7_datapath #(
      .ROWS(ROWS),
      .COLS(COLS)
  ) DATAPATH_7X7 (

      .clk(clk),
      .rst_n(rst_n),
      .d0_i(d0_i),
      .d1_i(d1_i),
      .d2_i(d2_i),
      .d3_i(d3_i),
      .d4_i(d4_i),
      .d5_i(d5_i),
      .d6_i(d6_i),
      .o_en(o_en),
      .d0_o(d0_o),
      .d1_o(d1_o),
      .d2_o(d2_o),
      .d3_o(d3_o),
      .d4_o(d4_o),
      .d5_o(d5_o),
      .d6_o(d6_o),
      .d7_o(d7_o),
      .d8_o(d8_o),
      .d9_o(d9_o),
      .d10_o(d10_o),
      .d11_o(d11_o),
      .d12_o(d12_o),
      .d13_o(d13_o),
      .d14_o(d14_o),
      .d15_o(d15_o),
      .d16_o(d16_o),
      .d17_o(d17_o),
      .d18_o(d18_o),
      .d19_o(d19_o),
      .d20_o(d20_o),
      .d21_o(d21_o),
      .d22_o(d22_o),
      .d23_o(d23_o),
      .d24_o(d24_o),
      .d25_o(d25_o),
      .d26_o(d26_o),
      .d27_o(d27_o),
      .d28_o(d28_o),
      .d29_o(d29_o),
      .d30_o(d30_o),
      .d31_o(d31_o),
      .d32_o(d32_o),
      .d33_o(d33_o),
      .d34_o(d34_o),
      .d35_o(d35_o),
      .d36_o(d36_o),
      .d37_o(d37_o),
      .d38_o(d38_o),
      .d39_o(d39_o),
      .d40_o(d40_o),
      .d41_o(d41_o),
      .d42_o(d42_o),
      .d43_o(d43_o),
      .d44_o(d44_o),
      .d45_o(d45_o),
      .d46_o(d46_o),
      .d47_o(d47_o),
      .d48_o(d48_o),
      .finish_en(finish_en),
      .padding_fi(padding_fi),
      .count_en(count_en),
      .reset_en(reset_en)
  );

endmodule
