module top_module #(
    parameter COLS = 128,
    parameter ROWS = 128
) (
    input clk,
    input rst_n,
    input start_i,
    // slave interface
    input [7:0] grayscale_i,
    input i_valid,
    output o_data_ready,
    // master interface 
    output [31:0] histogram_o,
    output o_valid,
    input i_data_ready,
    // interrupt
    output o_intr
);

  assign o_data_ready = 1'b1;

  wire axis_prog_full;

  wire finish;
  wire read_finish;
  wire read_en;
  wire [31:0] histogram;
  wire o_histogram_valid;
  wire o_intr_o;
  wire start_en;
  top_module__controller inst_top_module__controller (
      .clk        (clk),
      .rst_n      (rst_n),
      .finish_i   (finish),
      .start_en   (start_en),
      .read_finish(read_finish),
      .o_intr     (o_intr_o),
      .read_en    (read_en)
  );
  top_module__datapath #(
      .COLS(COLS),
      .ROWS(ROWS)
  ) inst_top_module__datapath (
      .clk        (clk),
      .rst_n      (rst_n),
      .grayscale_i(grayscale_i),
      .i_valid    (i_valid),
      .start_i    (start_i),
      .start_en   (start_en),
      .read_en    (read_en),
      .histogram_o(histogram),
      .o_valid    (o_histogram_valid),
      .finish     (finish),
      .read_finish(read_finish)
  );


  assign histogram_o = histogram;
  assign o_intr = o_intr_o;
  assign o_valid = o_histogram_valid;
  //   integer file;
  //   always @(posedge clk) begin
  //     if (~rst_n) begin
  //       file = $fopen("D:\\Thesis\\codetest\\python\\histogram_verilog_prev.txt", "w");
  //     end else if (o_histogram_valid) begin
  //       $fwrite(file, "%d\n", histogram);
  //     end else if (o_intr) begin
  //       $fclose(file);
  //     end
  //   end


endmodule

