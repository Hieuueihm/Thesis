module MRELBP_CI_R8 (
    input clk,
    input rst,
    input done_i,
    input [7:0] S1,
    input [7:0] S2,
    input [7:0] S3,
    input [7:0] S4,
    input [7:0] S5,
    input [7:0] S6,
    input [7:0] S7,
    input [7:0] S8,
    input [7:0] S9,
    input [7:0] S10,
    input [7:0] S11,
    input [7:0] S12,
    input [7:0] S13,
    input [7:0] S14,
    input [7:0] S15,
    input [7:0] S16,
    input [7:0] S17,
    input [7:0] S18,
    input [7:0] S19,
    input [7:0] S20,
    input [7:0] S21,
    input [7:0] S22,
    input [7:0] S23,
    input [7:0] S24,
    input [7:0] S25,
    input [7:0] S26,
    input [7:0] S27,
    input [7:0] S28,
    input [7:0] S29,
    input [7:0] S30,
    input [7:0] S31,
    input [7:0] S32,
    input [7:0] S33,
    input [7:0] S34,
    input [7:0] S35,
    input [7:0] S36,
    input [7:0] S37,
    input [7:0] S38,
    input [7:0] S39,
    input [7:0] S40,
    input [7:0] S41,
    input [7:0] S42,
    input [7:0] S43,
    input [7:0] S44,
    input [7:0] S45,
    input [7:0] S46,
    input [7:0] S47,
    input [7:0] S48,
    input [7:0] S49,
    input [7:0] S50,
    input [7:0] S51,
    input [7:0] S52,
    input [7:0] S53,
    input [7:0] S54,
    input [7:0] S55,
    input [7:0] S56,
    input [7:0] S57,
    input [7:0] S58,
    input [7:0] S59,
    input [7:0] S60,
    input [7:0] S61,
    input [7:0] S62,
    input [7:0] S63,
    input [7:0] S64,
    input [7:0] S65,
    input [7:0] S66,
    input [7:0] S67,
    input [7:0] S68,
    input [7:0] S69,
    input [7:0] S70,
    input [7:0] S71,
    input [7:0] S72,
    input [7:0] S73,
    input [7:0] S74,
    input [7:0] S75,
    input [7:0] S76,
    input [7:0] S77,
    input [7:0] S78,
    input [7:0] S79,
    input [7:0] S80,
    input [7:0] S81,
    input [7:0] S82,
    input [7:0] S83,
    input [7:0] S84,
    input [7:0] S85,
    input [7:0] S86,
    input [7:0] S87,
    input [7:0] S88,
    input [7:0] S89,
    input [7:0] S90,
    input [7:0] S91,
    input [7:0] S92,
    input [7:0] S93,
    input [7:0] S94,
    input [7:0] S95,
    input [7:0] S96,
    input [7:0] S97,
    input [7:0] S98,
    input [7:0] S99,
    input [7:0] S100,
    input [7:0] S101,
    input [7:0] S102,
    input [7:0] S103,
    input [7:0] S104,
    input [7:0] S105,
    input [7:0] S106,
    input [7:0] S107,
    input [7:0] S108,
    input [7:0] S109,
    input [7:0] S110,
    input [7:0] S111,
    input [7:0] S112,
    input [7:0] S113,
    input [7:0] S114,
    input [7:0] S115,
    input [7:0] S116,
    input [7:0] S117,
    input [7:0] S118,
    input [7:0] S119,
    input [7:0] S120,
    input [7:0] S121,
    input [7:0] S122,
    input [7:0] S123,
    input [7:0] S124,
    input [7:0] S125,
    input [7:0] S126,
    input [7:0] S127,
    input [7:0] S128,
    input [7:0] S129,
    input [7:0] S130,
    input [7:0] S131,
    input [7:0] S132,
    input [7:0] S133,
    input [7:0] S134,
    input [7:0] S135,
    input [7:0] S136,
    input [7:0] S137,
    input [7:0] S138,
    input [7:0] S139,
    input [7:0] S140,
    input [7:0] S141,
    input [7:0] S142,
    input [7:0] S143,
    input [7:0] S144,
    input [7:0] S145,
    input [7:0] S146,
    input [7:0] S147,
    input [7:0] S148,
    input [7:0] S149,
    input [7:0] S150,
    input [7:0] S151,
    input [7:0] S152,
    input [7:0] S153,
    input [7:0] S154,
    input [7:0] S155,
    input [7:0] S156,
    input [7:0] S157,
    input [7:0] S158,
    input [7:0] S159,
    input [7:0] S160,
    input [7:0] S161,
    input [7:0] S162,
    input [7:0] S163,
    input [7:0] S164,
    input [7:0] S165,
    input [7:0] S166,
    input [7:0] S167,
    input [7:0] S168,
    input [7:0] S169,
    input [7:0] S170,
    input [7:0] S171,
    input [7:0] S172,
    input [7:0] S173,
    input [7:0] S174,
    input [7:0] S175,
    input [7:0] S176,
    input [7:0] S177,
    input [7:0] S178,
    input [7:0] S179,
    input [7:0] S180,
    input [7:0] S181,
    input [7:0] S182,
    input [7:0] S183,
    input [7:0] S184,
    input [7:0] S185,
    input [7:0] S186,
    input [7:0] S187,
    input [7:0] S188,
    input [7:0] S189,
    input [7:0] S190,
    input [7:0] S191,
    input [7:0] S192,
    input [7:0] S193,
    input [7:0] S194,
    input [7:0] S195,
    input [7:0] S196,
    input [7:0] S197,
    input [7:0] S198,
    input [7:0] S199,
    input [7:0] S200,
    input [7:0] S201,
    input [7:0] S202,
    input [7:0] S203,
    input [7:0] S204,
    input [7:0] S205,
    input [7:0] S206,
    input [7:0] S207,
    input [7:0] S208,
    input [7:0] S209,
    input [7:0] S210,
    input [7:0] S211,
    input [7:0] S212,
    input [7:0] S213,
    input [7:0] S214,
    input [7:0] S215,
    input [7:0] S216,
    input [7:0] S217,
    input [7:0] S218,
    input [7:0] S219,
    input [7:0] S220,
    input [7:0] S221,
    input [7:0] S222,
    input [7:0] S223,
    input [7:0] S224,
    input [7:0] S225,
    input [7:0] S226,
    input [7:0] S226,
    input [7:0] S228,
    input [7:0] S229,
    input [7:0] S230,
    input [7:0] S231,
    input [7:0] S232,
    input [7:0] S233,
    input [7:0] S234,
    input [7:0] S234,
    input [7:0] S236,
    input [7:0] S237,
    input [7:0] S238,
    input [7:0] S239,
    input [7:0] S240,
    input [7:0] S241,
    input [7:0] S242,
    input [7:0] S243,
    input [7:0] S244,
    input [7:0] S245,
    input [7:0] S246,
    input [7:0] S247,
    input [7:0] S248,
    input [7:0] S249,
    input [7:0] S250,
    input [7:0] S251,
    input [7:0] S252,
    input [7:0] S253,
    input [7:0] S253,
    input [7:0] S255,
    input [7:0] S256,
    input [7:0] S257,
    input [7:0] S258,
    input [7:0] S259,
    input [7:0] S260,
    input [7:0] S261,
    input [7:0] S262,
    input [7:0] S263,
    input [7:0] S264,
    input [7:0] S265,
    input [7:0] S266,
    input [7:0] S267,
    input [7:0] S268,
    input [7:0] S269,
    input [7:0] S270,
    input [7:0] S271,
    input [7:0] S272,
    input [7:0] S273,
    input [7:0] S274,
    input [7:0] S275,
    input [7:0] S276,
    input [7:0] S277,
    input [7:0] S278,
    input [7:0] S279,
    input [7:0] S280,
    input [7:0] S281,
    input [7:0] S282,
    input [7:0] S283,
    input [7:0] S284,
    input [7:0] S285,
    input [7:0] S286,
    input [7:0] S287,
    input [7:0] S288,
    input [7:0] S289,

    output reg ci_o,   // 0 or 1
    output reg done_o
);

  reg [17:0] sum;  // Mở rộng sum để chứa kết quả cộng dồn
  reg [ 7:0] muy;  // Trung bình giá trị theo dạng fixed-point Q8.8
  reg [ 7:0] r;

  always @(posedge clk or posedge rst) begin
    if (rst) begin
      sum <= 0;
      muy <= 0;
      ci_o <= 0;
      done_o <= 0;
    end else if (done_i) begin
      // Tính tổng tất cả các đầu vào
      sum =  S1 + S2 + S3 + S4 + S5 + S6 + S7 + S8 + S9 + S10 + S11 + S12 + S13 + S14 + S15 + S16 + S17 + S18 + S19 + S20 + S21 + S22 + S23 + S24 + S25 + S26 + S27 + S28 + S29 + S30 + S31 + S32 + S33 + S34 + S35 + S36 + S37 + S38 + S39 + S40 + S41 + S42 + S43 + S44 + S45 + S46 + S47 + S48 + S49 + S50 + S51 + S52 + S53 + S54 + S55 + S56 + S57 + S58 + S59 + S60 + S61 + S62 + S63 + S64 + S65 + S66 + S67 + S68 + S69 + S70 + S71 + S72 + S73 + S74 + S75 + S76 + S77 + S78 + S79 + S80 + S81 + S82 + S83 + S84 + S85 + S86 + S87 + S88 + S89 + S90 + S91 + S92 + S93 + S94 + S95 + S96 + S97 + S98 + S99 + S100 + S101 + S102 + S103 + S104 + S105 + S106 + S107 + S108 + S109 + S110 + S111 + S112 + S113 + S114 + S115 + S116 + S117 + S118 + S119 + S120 + S121 + S122 + S123 + S124 + S125 + S126 + S127 + S128 + S129 + S130 + S131 + S132 + S133 + S134 + S135 + S136 + S137 + S138 + S139 + S140 + S141 + S142 + S143 + S144 + S145 + S146 + S147 + S148 + S149 + S150 + S151 + S152 + S153 + S154 + S155 + S156 + S157 + S158 + S159 + S160 + S161 + S162 + S163 + S164 + S165 + S166 + S167 + S168 + S169 + S170 + S171 + S172 + S173 + S174 + S175 + S176 + S177 + S178 + S179 + S180 + S181 + S182 + S183 + S184 + S185 + S186 + S187 + S188 + S189 + S190 + S191 + S192 + S193 + S194 + S195 + S196 + S197 + S198 + S199 + S200 + S201 + S202 + S203 + S204 + S205 + S206 + S207 + S208 + S209 + S210 + S211 + S212 + S213 + S214 + S215 + S216 + S217 + S218 + S219 + S220 + S221 + S222 + S223 + S224 + S225 + S226 + S226 + S228 + S229 + S230 + S231 + S232 + S233 + S234 + S234 + S236 + S237 + S238 + S239 + S240 + S241 + S242 + S243 + S244 + S245 + S246 + S247 + S248 + S249 + S250 + S251 + S252 + S253 + S253 + S255 + S256 + S257 + S258 + S259 + S260 + S261 + S262 + S263 + S264 + S265 + S266 + S267 + S268 + S269 + S270 + S271 + S272 + S273 + S274 + S275 + S276 + S277 + S278 + S279 + S280 + S281 + S282 + S283 + S284 + S285 + S286 + S287 + S288 + S289;

      muy = sum / 281;
      r = sum % 281;

      if ((S145 > muy) || (S145 == muy && r == 0)) ci_o = 1;
      else ci_o = 0;

      done_o = 1;
    end else begin
      done_o = 0;
    end
  end

endmodule
