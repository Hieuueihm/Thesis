function int get_template_id();
// Template 0 - Center (0,0)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o == 0 &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o == 0 &&
    vif.d11_o == 0 &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 0;
// Template 1 - Center (0,1)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o == 0 &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o == 0 &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 1;
// Template 2 - Center (0,2)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o == 0 &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 2;
// Template 3 - Center (0,5)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o == 0 &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o == 0
) return 3;
// Template 4 - Center (0,6)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o == 0 &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o == 0 &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 4;
// Template 5 - Center (1,0)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o == 0 &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 5;
// Template 6 - Center (1,1)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o == 0 &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 6;
// Template 7 - Center (1,2)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 7;
// Template 8 - Center (1,5)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o == 0
) return 8;
// Template 9 - Center (1,6)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o == 0 &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o == 0 &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 9;
// Template 10 - Center (2,0)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o == 0 &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 10;
// Template 11 - Center (2,1)
if (
    vif.d0_o == 0 &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 11;
// Template 12 - Center (2,2)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o inside {[0:255]}
) return 12;
// Template 13 - Center (2,5)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o inside {[0:255]} &&
    vif.d24_o == 0
) return 13;
// Template 14 - Center (2,6)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o == 0 &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o inside {[0:255]} &&
    vif.d21_o inside {[0:255]} &&
    vif.d22_o inside {[0:255]} &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 14;
// Template 15 - Center (5,0)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o == 0 &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 15;
// Template 16 - Center (5,1)
if (
    vif.d0_o == 0 &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 16;
// Template 17 - Center (5,2)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o inside {[0:255]} &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 17;
// Template 18 - Center (5,5)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o inside {[0:255]} &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 18;
// Template 19 - Center (5,6)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o == 0 &&
    vif.d14_o == 0 &&
    vif.d15_o inside {[0:255]} &&
    vif.d16_o inside {[0:255]} &&
    vif.d17_o inside {[0:255]} &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 19;
// Template 20 - Center (6,0)
if (
    vif.d0_o == 0 &&
    vif.d1_o == 0 &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o == 0 &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o == 0 &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o == 0 &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 20;
// Template 21 - Center (6,1)
if (
    vif.d0_o == 0 &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o == 0 &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o == 0 &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o == 0 &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 21;
// Template 22 - Center (6,2)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o inside {[0:255]} &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o inside {[0:255]} &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o inside {[0:255]} &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o == 0 &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 22;
// Template 23 - Center (6,5)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o inside {[0:255]} &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o inside {[0:255]} &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o inside {[0:255]} &&
    vif.d14_o == 0 &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o == 0 &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 23;
// Template 24 - Center (6,6)
if (
    vif.d0_o inside {[0:255]} &&
    vif.d1_o inside {[0:255]} &&
    vif.d2_o inside {[0:255]} &&
    vif.d3_o == 0 &&
    vif.d4_o == 0 &&
    vif.d5_o inside {[0:255]} &&
    vif.d6_o inside {[0:255]} &&
    vif.d7_o inside {[0:255]} &&
    vif.d8_o == 0 &&
    vif.d9_o == 0 &&
    vif.d10_o inside {[0:255]} &&
    vif.d11_o inside {[0:255]} &&
    vif.d12_o inside {[0:255]} &&
    vif.d13_o == 0 &&
    vif.d14_o == 0 &&
    vif.d15_o == 0 &&
    vif.d16_o == 0 &&
    vif.d17_o == 0 &&
    vif.d18_o == 0 &&
    vif.d19_o == 0 &&
    vif.d20_o == 0 &&
    vif.d21_o == 0 &&
    vif.d22_o == 0 &&
    vif.d23_o == 0 &&
    vif.d24_o == 0
) return 24;
else return -1;
endfunction