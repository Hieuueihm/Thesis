`timescale 1ns / 1ps

module sum_cumulative_top_tb();
    reg clk; reg rst; reg done_i;
    reg [9:0] i_col;
    reg [7:0] S1, S2, S3, S4, S5, S6, S7, S8, S9, S10;
    reg [7:0] S11, S12, S13, S14, S15, S16, S17, S18, S19, S20; reg [7:0] S21, S22, S23, S24, S25;
    wire [12:0] sum_o;
    wire done_o;
    sum_cumulative_top uut
    (.clk(clk), .rst(rst), .done_i(done_i), .i_col(i_col), .S1(S1), .S2(S2), .S3(S3), .S4(S4), .S5(S5), .S6(S6), .S7(S7), .S8(S8), .S9(S9),
    .S10(S10), .S11(S11), .S12(S12), .S13(S13), .S14(S14), .S15(S15), .S16(S16), .S17(S17), .S18(S18), .S19(S19), .S20(S20), .S21(S21), .S22(S22),
    .S23(S23), .S24(S24), .S25(S25), .sum_o(sum_o),.done_o(done_o));
    
    // Clock generation
    initial clk   = 0;
    always #5 clk = ~clk; // 100MHz clock
    
    // Test stimulus
    initial begin
        // Initialize inputs
        rst    = 1;
        done_i = 0;
        S1     = 8'd0; S2     = 8'd0; S3     = 8'd0; S4     = 8'd0; S5     = 8'd0;
        S6     = 8'd0; S7     = 8'd0; S8     = 8'd0; S9     = 8'd0; S10     = 8'd0;
        S11    = 8'd0; S12    = 8'd0; S13    = 8'd0; S14    = 8'd0; S15    = 8'd0;
        S16    = 8'd0; S17    = 8'd0; S18    = 8'd0; S19    = 8'd0; S20    = 8'd0;
        S21    = 8'd0; S22    = 8'd0; S23    = 8'd0; S24    = 8'd0; S25    = 8'd0;
        
        // Apply reset
        #10 rst = 0;
        
        // Apply stimulus
        #10 done_i = 1;
        i_col      = 10'd0;
        S1         = 8'd1; S2         = 8'd2; S3         = 8'd3; S4         = 8'd4; S5         = 8'd5;
        S6         = 8'd6; S7         = 8'd7; S8         = 8'd8; S9         = 8'd9; S10         = 8'd10;
        S11        = 8'd11; S12        = 8'd12; S13        = 8'd13; S14        = 8'd14; S15        = 8'd15;
        S16        = 8'd16; S17        = 8'd17; S18        = 8'd18; S19        = 8'd19; S20        = 8'd20;
        S21        = 8'd21; S22        = 8'd22; S23        = 8'd23; S24        = 8'd24; S25        = 8'd25;
        
        // sum = 325
        
        #10;
        i_col = 10'd1;
        S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd12;
        S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd13;
        S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd14;
        S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd100;
        S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd200;
        #10;
        i_col = 10'd2;
        S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd15;
        S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd15;
        S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd15;
        S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd15;
        S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd0;
        #10;
        i_col = 10'd2;
        S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd100;
        S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd100;
        S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd100;
        S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd100;
        S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd0;
        #10;
        i_col = 10'd0;
        S1    = 8'd10; S2    = 8'd10; S3    = 8'd10; S4    = 8'd10; S5    = 8'd10;
        S6    = 8'd10; S7    = 8'd10; S8    = 8'd10; S9    = 8'd10; S10    = 8'd10;
        S11   = 8'd10; S12   = 8'd10; S13   = 8'd10; S14   = 8'd10; S15   = 8'd10;
        S16   = 8'd10; S17   = 8'd10; S18   = 8'd10; S19   = 8'd10; S20   = 8'd10;
        S21   = 8'd10; S22   = 8'd10; S23   = 8'd10; S24   = 8'd10; S25   = 8'd10;
        #10;
        i_col = 10'd1;
        S1    = 8'd10; S2    = 8'd10; S3    = 8'd10; S4    = 8'd10; S5    = 8'd20;
        S6    = 8'd10; S7    = 8'd10; S8    = 8'd10; S9    = 8'd10; S10    = 8'd20;
        S11   = 8'd10; S12   = 8'd10; S13   = 8'd10; S14   = 8'd10; S15   = 8'd20;
        S16   = 8'd10; S17   = 8'd10; S18   = 8'd10; S19   = 8'd10; S20   = 8'd20;
        S21   = 8'd10; S22   = 8'd10; S23   = 8'd10; S24   = 8'd10; S25   = 8'd20;
        #10;
        done_i = 0;
        // // Wait for some cycles
        // #10;
        // i_col = 10'd2;
        // S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd3;
        // S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd11;
        // S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd14;
        // S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd10;
        // S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd200;
        // #10;
        // i_col = 10'd3;
        // S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd14;
        // S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd3;
        // S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd19;
        // S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd10;
        // S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd20;
        // #10;
        // i_col = 10'd4;
        // S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd12;
        // S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd13;
        // S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd16;
        // S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd18;
        // S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd22;
        // #10;
        // i_col = 10'd0;
        // S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd19;
        // S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd21;
        // S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd22;
        // S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd32;
        // S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd33;
        // #10;
        // i_col = 10'd1;
        // S1    = 8'd1; S2    = 8'd2; S3    = 8'd3; S4    = 8'd4; S5    = 8'd22;
        // S6    = 8'd6; S7    = 8'd7; S8    = 8'd8; S9    = 8'd9; S10    = 8'd26;
        // S11   = 8'd11; S12   = 8'd12; S13   = 8'd13; S14   = 8'd14; S15   = 8'd22;
        // S16   = 8'd16; S17   = 8'd17; S18   = 8'd18; S19   = 8'd19; S20   = 8'd32;
        // S21   = 8'd21; S22   = 8'd22; S23   = 8'd23; S24   = 8'd24; S25   = 8'd33;
        #200;
        
        
        
        // Add more stimulus if needed
        
        // Finish simulation
        #100 $stop;
    end
    
endmodule
