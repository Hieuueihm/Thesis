// R = 2 ->  (2* 2 + 1)^2 = 25
module MRELBP_CI_R2 (
    input clk,
    input rst,
    input done_i,
    input [7:0] S1,
    input [7:0] S2,
    input [7:0] S3,
    input [7:0] S4,
    input [7:0] S5,
    input [7:0] S6,
    input [7:0] S7,
    input [7:0] S8,
    input [7:0] S9,
    output [7:0] ci_o,
    output reg done_o
);  // 255 * 8 = 

  function [0:0] sign_function(input signed [8:0] input_value);
    begin
      if (input_value >= 0) begin
        sign_function = 1'b1;
      end else begin
        sign_function = 1'b0;
      end
    end
  endfunction
  reg [10:0] sum;
  reg [ 8:0] muy;
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      ci_o   <= 8'b0;
      done_o <= 0;
    end else if (done_i) begin
      sum = S1 + S2 + S3 + S4 + S5 + S6 + S7 + S8 + S9;

      // muy = (sum >> 4) + (sum >> 5) + (sum >> 6);  // optimize after
      muy = sum / 9;
      ci_o = sign_function(S5 - muy);
      done_o = 1;
    end else begin
      done_o <= 0;
    end
  end



endmodule
