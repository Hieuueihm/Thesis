module Window_buffer_15x15 #(parameter COLS = 11,
                             parameter ROWS = 11)
                            (input clk,
                             input rst,
                             input done_i,
                             input[7:0] S1_i,
                             S2_i,
                             S3_i,
                             S4_i,
                             S5_i,
                             S6_i,
                             S7_i,
                             S8_i,
                             S9_i,
                             S10_i,
                             S11_i,
                             S12_i,
                             S13_i,
                             S14_i,
                             S15_i,
                             output[7:0] S1_o,
                             S2_o,
                             S3_o,
                             S4_o,
                             S5_o,
                             S6_o,
                             S7_o,
                             S8_o,
                             S9_o,
                             S10_o,
                             S11_o,
                             S12_o,
                             S13_o,
                             S14_o,
                             S15_o,
                             S16_o,
                             S17_o,
                             S18_o,
                             S19_o,
                             S20_o,
                             S21_o,
                             S22_o,
                             S23_o,
                             S24_o,
                             S25_o,
                             S26_o,
                             S27_o,
                             S28_o,
                             S29_o,
                             S30_o,
                             S31_o,
                             S32_o,
                             S33_o,
                             S34_o,
                             S35_o,
                             S36_o,
                             S37_o,
                             S38_o,
                             S39_o,
                             S40_o,
                             S41_o,
                             S42_o,
                             S43_o,
                             S44_o,
                             S45_o,
                             S46_o,
                             S47_o,
                             S48_o,
                             S49_o,
                             S50_o,
                             S51_o,
                             S52_o,
                             S53_o,
                             S54_o,
                             S55_o,
                             S56_o,
                             S57_o,
                             S58_o,
                             S59_o,
                             S60_o,
                             S61_o,
                             S62_o,
                             S63_o,
                             S64_o,
                             S65_o,
                             S66_o,
                             S67_o,
                             S68_o,
                             S69_o,
                             S70_o,
                             S71_o,
                             S72_o,
                             S73_o,
                             S74_o,
                             S75_o,
                             S76_o,
                             S77_o,
                             S78_o,
                             S79_o,
                             S80_o,
                             S81_o,
                             S82_o,
                             S83_o,
                             S84_o,
                             S85_o,
                             S86_o,
                             S87_o,
                             S88_o,
                             S89_o,
                             S90_o,
                             S91_o,
                             S92_o,
                             S93_o,
                             S94_o,
                             S95_o,
                             S96_o,
                             S97_o,
                             S98_o,
                             S99_o,
                             S100_o,
                             S101_o,
                             S102_o,
                             S103_o,
                             S104_o,
                             S105_o,
                             S106_o,
                             S107_o,
                             S108_o,
                             S109_o,
                             S110_o,
                             S111_o,
                             S112_o,
                             S113_o,
                             S114_o,
                             S115_o,
                             S116_o,
                             S117_o,
                             S118_o,
                             S119_o,
                             S120_o,
                             S121_o,
                             S122_o,
                             S123_o,
                             S124_o,
                             S125_o,
                             S126_o,
                             S127_o,
                             S128_o,
                             S129_o,
                             S130_o,
                             S131_o,
                             S132_o,
                             S133_o,
                             S134_o,
                             S135_o,
                             S136_o,
                             S137_o,
                             S138_o,
                             S139_o,
                             S140_o,
                             S141_o,
                             S142_o,
                             S143_o,
                             S144_o,
                             S145_o,
                             S146_o,
                             S147_o,
                             S148_o,
                             S149_o,
                             S150_o,
                             S151_o,
                             S152_o,
                             S153_o,
                             S154_o,
                             S155_o,
                             S156_o,
                             S157_o,
                             S158_o,
                             S159_o,
                             S160_o,
                             S161_o,
                             S162_o,
                             S163_o,
                             S164_o,
                             S165_o,
                             S166_o,
                             S167_o,
                             S168_o,
                             S169_o,
                             S170_o,
                             S171_o,
                             S172_o,
                             S173_o,
                             S174_o,
                             S175_o,
                             S176_o,
                             S177_o,
                             S178_o,
                             S179_o,
                             S180_o,
                             S181_o,
                             S182_o,
                             S183_o,
                             S184_o,
                             S185_o,
                             S186_o,
                             S187_o,
                             S188_o,
                             S189_o,
                             S190_o,
                             S191_o,
                             S192_o,
                             S193_o,
                             S194_o,
                             S195_o,
                             S196_o,
                             S197_o,
                             S198_o,
                             S199_o,
                             S200_o,
                             S201_o,
                             S202_o,
                             S203_o,
                             S204_o,
                             S205_o,
                             S206_o,
                             S207_o,
                             S208_o,
                             S209_o,
                             S210_o,
                             S211_o,
                             S212_o,
                             S213_o,
                             S214_o,
                             S215_o,
                             S216_o,
                             S217_o,
                             S218_o,
                             S219_o,
                             S220_o,
                             S221_o,
                             S222_o,
                             S223_o,
                             S224_o,
                             S225_o,
                             output done_o,
                             output progress_done_o);
    wire i_row_eq_max, i_col_eq_max, i_col_ge_threshold;
    wire count_en;
    
    Window_buffer_15x15_datapath #(
    .COLS(COLS),
    .ROWS(ROWS)
    ) inst_Window_buffer_15x15_datapath (
    .clk                (clk),
    .rst                (rst),
    .count_en           (count_en),
    .S1_i               (S1_i),
    .S2_i               (S2_i),
    .S3_i               (S3_i),
    .S4_i               (S4_i),
    .S5_i               (S5_i),
    .S6_i               (S6_i),
    .S7_i               (S7_i),
    .S8_i               (S8_i),
    .S9_i               (S9_i),
    .S10_i              (S10_i),
    .S11_i              (S11_i),
    .S12_i              (S12_i),
    .S13_i              (S13_i),
    .S14_i              (S14_i),
    .S15_i              (S15_i),
    .i_row_eq_max       (i_row_eq_max),
    .S1_o               (S1_o),
    .S2_o               (S2_o),
    .S3_o               (S3_o),
    .S4_o               (S4_o),
    .S5_o               (S5_o),
    .S6_o               (S6_o),
    .S7_o               (S7_o),
    .S8_o               (S8_o),
    .S9_o               (S9_o),
    .S10_o              (S10_o),
    .S11_o              (S11_o),
    .S12_o              (S12_o),
    .S13_o              (S13_o),
    .S14_o              (S14_o),
    .S15_o              (S15_o),
    .S16_o              (S16_o),
    .S17_o              (S17_o),
    .S18_o              (S18_o),
    .S19_o              (S19_o),
    .S20_o              (S20_o),
    .S21_o              (S21_o),
    .S22_o              (S22_o),
    .S23_o              (S23_o),
    .S24_o              (S24_o),
    .S25_o              (S25_o),
    .S26_o              (S26_o),
    .S27_o              (S27_o),
    .S28_o              (S28_o),
    .S29_o              (S29_o),
    .S30_o              (S30_o),
    .S31_o              (S31_o),
    .S32_o              (S32_o),
    .S33_o              (S33_o),
    .S34_o              (S34_o),
    .S35_o              (S35_o),
    .S36_o              (S36_o),
    .S37_o              (S37_o),
    .S38_o              (S38_o),
    .S39_o              (S39_o),
    .S40_o              (S40_o),
    .S41_o              (S41_o),
    .S42_o              (S42_o),
    .S43_o              (S43_o),
    .S44_o              (S44_o),
    .S45_o              (S45_o),
    .S46_o              (S46_o),
    .S47_o              (S47_o),
    .S48_o              (S48_o),
    .S49_o              (S49_o),
    .S50_o              (S50_o),
    .S51_o              (S51_o),
    .S52_o              (S52_o),
    .S53_o              (S53_o),
    .S54_o              (S54_o),
    .S55_o              (S55_o),
    .S56_o              (S56_o),
    .S57_o              (S57_o),
    .S58_o              (S58_o),
    .S59_o              (S59_o),
    .S60_o              (S60_o),
    .S61_o              (S61_o),
    .S62_o              (S62_o),
    .S63_o              (S63_o),
    .S64_o              (S64_o),
    .S65_o              (S65_o),
    .S66_o              (S66_o),
    .S67_o              (S67_o),
    .S68_o              (S68_o),
    .S69_o              (S69_o),
    .S70_o              (S70_o),
    .S71_o              (S71_o),
    .S72_o              (S72_o),
    .S73_o              (S73_o),
    .S74_o              (S74_o),
    .S75_o              (S75_o),
    .S76_o              (S76_o),
    .S77_o              (S77_o),
    .S78_o              (S78_o),
    .S79_o              (S79_o),
    .S80_o              (S80_o),
    .S81_o              (S81_o),
    .S82_o              (S82_o),
    .S83_o              (S83_o),
    .S84_o              (S84_o),
    .S85_o              (S85_o),
    .S86_o              (S86_o),
    .S87_o              (S87_o),
    .S88_o              (S88_o),
    .S89_o              (S89_o),
    .S90_o              (S90_o),
    .S91_o              (S91_o),
    .S92_o              (S92_o),
    .S93_o              (S93_o),
    .S94_o              (S94_o),
    .S95_o              (S95_o),
    .S96_o              (S96_o),
    .S97_o              (S97_o),
    .S98_o              (S98_o),
    .S99_o              (S99_o),
    .S100_o             (S100_o),
    .S101_o             (S101_o),
    .S102_o             (S102_o),
    .S103_o             (S103_o),
    .S104_o             (S104_o),
    .S105_o             (S105_o),
    .S106_o             (S106_o),
    .S107_o             (S107_o),
    .S108_o             (S108_o),
    .S109_o             (S109_o),
    .S110_o             (S110_o),
    .S111_o             (S111_o),
    .S112_o             (S112_o),
    .S113_o             (S113_o),
    .S114_o             (S114_o),
    .S115_o             (S115_o),
    .S116_o             (S116_o),
    .S117_o             (S117_o),
    .S118_o             (S118_o),
    .S119_o             (S119_o),
    .S120_o             (S120_o),
    .S121_o             (S121_o),
    .S122_o             (S122_o),
    .S123_o             (S123_o),
    .S124_o             (S124_o),
    .S125_o             (S125_o),
    .S126_o             (S126_o),
    .S127_o             (S127_o),
    .S128_o             (S128_o),
    .S129_o             (S129_o),
    .S130_o             (S130_o),
    .S131_o             (S131_o),
    .S132_o             (S132_o),
    .S133_o             (S133_o),
    .S134_o             (S134_o),
    .S135_o             (S135_o),
    .S136_o             (S136_o),
    .S137_o             (S137_o),
    .S138_o             (S138_o),
    .S139_o             (S139_o),
    .S140_o             (S140_o),
    .S141_o             (S141_o),
    .S142_o             (S142_o),
    .S143_o             (S143_o),
    .S144_o             (S144_o),
    .S145_o             (S145_o),
    .S146_o             (S146_o),
    .S147_o             (S147_o),
    .S148_o             (S148_o),
    .S149_o             (S149_o),
    .S150_o             (S150_o),
    .S151_o             (S151_o),
    .S152_o             (S152_o),
    .S153_o             (S153_o),
    .S154_o             (S154_o),
    .S155_o             (S155_o),
    .S156_o             (S156_o),
    .S157_o             (S157_o),
    .S158_o             (S158_o),
    .S159_o             (S159_o),
    .S160_o             (S160_o),
    .S161_o             (S161_o),
    .S162_o             (S162_o),
    .S163_o             (S163_o),
    .S164_o             (S164_o),
    .S165_o             (S165_o),
    .S166_o             (S166_o),
    .S167_o             (S167_o),
    .S168_o             (S168_o),
    .S169_o             (S169_o),
    .S170_o             (S170_o),
    .S171_o             (S171_o),
    .S172_o             (S172_o),
    .S173_o             (S173_o),
    .S174_o             (S174_o),
    .S175_o             (S175_o),
    .S176_o             (S176_o),
    .S177_o             (S177_o),
    .S178_o             (S178_o),
    .S179_o             (S179_o),
    .S180_o             (S180_o),
    .S181_o             (S181_o),
    .S182_o             (S182_o),
    .S183_o             (S183_o),
    .S184_o             (S184_o),
    .S185_o             (S185_o),
    .S186_o             (S186_o),
    .S187_o             (S187_o),
    .S188_o             (S188_o),
    .S189_o             (S189_o),
    .S190_o             (S190_o),
    .S191_o             (S191_o),
    .S192_o             (S192_o),
    .S193_o             (S193_o),
    .S194_o             (S194_o),
    .S195_o             (S195_o),
    .S196_o             (S196_o),
    .S197_o             (S197_o),
    .S198_o             (S198_o),
    .S199_o             (S199_o),
    .S200_o             (S200_o),
    .S201_o             (S201_o),
    .S202_o             (S202_o),
    .S203_o             (S203_o),
    .S204_o             (S204_o),
    .S205_o             (S205_o),
    .S206_o             (S206_o),
    .S207_o             (S207_o),
    .S208_o             (S208_o),
    .S209_o             (S209_o),
    .S210_o             (S210_o),
    .S211_o             (S211_o),
    .S212_o             (S212_o),
    .S213_o             (S213_o),
    .S214_o             (S214_o),
    .S215_o             (S215_o),
    .S216_o             (S216_o),
    .S217_o             (S217_o),
    .S218_o             (S218_o),
    .S219_o             (S219_o),
    .S220_o             (S220_o),
    .S221_o             (S221_o),
    .S222_o             (S222_o),
    .S223_o             (S223_o),
    .S224_o             (S224_o),
    .S225_o             (S225_o),
    .i_col_eq_max       (i_col_eq_max),
    .i_col_ge_threshold (i_col_ge_threshold)
    );
    
    
    Window_buffer_15x15_controller inst_Window_buffer_15x15_controller (
    .clk                (clk),
    .rst                (rst),
    .done_i             (done_i),
    .i_row_eq_max       (i_row_eq_max),
    .i_col_eq_max       (i_col_eq_max),
    .i_col_ge_threshold (i_col_ge_threshold),
    .count_en           (count_en),
    .progress_done      (progress_done_o),
    .done_o             (done_o)
    );
    
    
endmodule
