module test(input clk,
            input rst,
            input [7:0] grayscale_i,
            input done_i);
    
    wire done_original_o;
    wire [7:0] data_o;
    wire done_3x3_o;
    wire [7:0] m_3x3_o;
    
    Median_processing #(.ROWS(30), .COLS(30))
    MEDIAN_PROCESSING
    (
    .clk(clk),
    .rst(rst),
    .data_i(grayscale_i),
    .done_i(done_i),
    .data_o(data_o),
    .done_o(done_original_o),
    .m_3x3_o(m_3x3_o),
    .done_3x3_o(done_3x3_o),
    .m_5x5_o(),
    .done_5x5_o(),
    .m_7x7_o(),
    .done_7x7_o(),
    .m_9x9_o(),
    .done_9x9_o()
    );
    
    wire [7:0] data0_3x3_o, data1_3x3_o, data2_3x3_o, data3_3x3_o, data4_3x3_o;
    wire done_buffer_3x3_o;
    Buffer_4_rows #(.DEPTH(30)) BUFFER_4_ROWS_3X3 (
    .clk(clk),
    .rst(rst),
    .done_i(done_3x3_o),
    .data_i(m_3x3_o),
    .data0_o(data0_3x3_o),
    .data1_o(data1_3x3_o),
    .data2_o(data2_3x3_o),
    .data3_o(data3_3x3_o),
    .data4_o(data4_3x3_o),
    .done_o(done_buffer_3x3_o)
    );
    
    wire [7:0] data0_o, data1_o, data2_o, data3_o, data4_o;
    wire done_o;
    Buffer_4_rows #(.DEPTH(30)) BUFFER_4_ROWS (
    .clk(clk),
    .rst(rst),
    .done_i(done_original_o),
    .data_i(data_o),
    .data0_o(data0_o),
    .data1_o(data1_o),
    .data2_o(data2_o),
    .data3_o(data3_o),
    .data4_o(data4_o),
    .done_o(done_o)
    );
    
    wire [7:0] data0_delay, data1_delay, data2_delay, data3_delay, data4_delay;
    shift_registers #(.WIDTH(8), .CYCLE(6))
    SHIFT_5_DATA0 (
    .clk(clk),
    .rst(rst),
    .data_i(data0_o),
    .data_o(data0_delay)
    );
    
    shift_registers #(.WIDTH(8), .CYCLE(6))
    SHIFT_5_DATA1 (
    .clk(clk),
    .rst(rst),
    .data_i(data1_o),
    .data_o(data1_delay)
    );
    
    
    shift_registers #(.WIDTH(8), .CYCLE(6))
    SHIFT_5_DATA2 (
    .clk(clk),
    .rst(rst),
    .data_i(data2_o),
    .data_o(data2_delay)
    );
    
    
    shift_registers #(.WIDTH(8), .CYCLE(6))
    SHIFT_5_DATA3 (
    .clk(clk),
    .rst(rst),
    .data_i(data3_o),
    .data_o(data3_delay)
    );
    
    shift_registers #(.WIDTH(8), .CYCLE(6))
    SHIFT_5_DATA4 (
    .clk(clk),
    .rst(rst),
    .data_i(data4_o),
    .data_o(data4_delay)
    );
    
    
    
endmodule
