module MRELBP_CI_R2_datapath (
    input clk,
    input rst,
    input s_all_en,
    input accum_en,
    input [7:0] data0_i,
    data1_i,
    data2_i,
    data3_i,
    data4_i,
    output reg ci_o,
    output reg done_o
);
  reg [7:0] p1_d0, p1_d1, p1_d2, p1_d3, p1_d4;
  reg [7:0] p2_d0, p2_d1, p2_d2, p2_d3, p2_d4;
  reg [7:0] p3_d0, p3_d1, p3_d2, p3_d3, p3_d4;
  reg [7:0] p4_d0, p4_d1, p4_d2, p4_d3, p4_d4;
  reg [7:0] p5_d0, p5_d1, p5_d2, p5_d3, p5_d4;

  reg [10:0] sum1, sum2, sum3, sum4, sum5;

  assign sum1 = (p1_d0 + p1_d1 + p1_d2 + p1_d3 + p1_d4);
  assign sum2 = (p2_d0 + p2_d1 + p2_d2 + p2_d3 + p2_d4);
  assign sum3 = (p3_d0 + p3_d1 + p3_d2 + p3_d3 + p3_d4);
  assign sum4 = (p4_d0 + p4_d1 + p4_d2 + p4_d3 + p4_d4);
  assign sum5 = (p5_d0 + p5_d1 + p5_d2 + p5_d3 + p5_d4);

  reg [15:0] sum_a;
  reg [15:0] muy;


  always @(posedge clk) begin
    if (rst) begin

      p1_d0  <= 0;
      p1_d1  <= 0;
      p1_d2  <= 0;
      p1_d3  <= 0;
      p1_d4  <= 0;

      p2_d0  <= 0;
      p2_d1  <= 0;
      p2_d2  <= 0;
      p2_d3  <= 0;
      p2_d4  <= 0;

      p3_d0  <= 0;
      p3_d1  <= 0;
      p3_d2  <= 0;
      p3_d3  <= 0;
      p3_d4  <= 0;

      p4_d0  <= 0;
      p4_d1  <= 0;
      p4_d2  <= 0;
      p4_d3  <= 0;
      p4_d4  <= 0;

      p5_d0  <= 0;
      p5_d1  <= 0;
      p5_d2  <= 0;
      p5_d3  <= 0;
      p5_d4  <= 0;

      ci_o   <= 0;
      done_o <= 0;
    end else begin
      p1_d0 <= data0_i;
      p1_d1 <= data1_i;
      p1_d2 <= data2_i;
      p1_d3 <= data3_i;
      p1_d4 <= data4_i;

      p2_d0 <= p1_d0;
      p2_d1 <= p1_d1;
      p2_d2 <= p1_d2;
      p2_d3 <= p1_d3;
      p2_d4 <= p1_d4;


      p3_d0 <= p2_d0;
      p3_d1 <= p2_d1;
      p3_d2 <= p2_d2;
      p3_d3 <= p2_d3;
      p3_d4 <= p2_d4;

      p4_d0 <= p3_d0;
      p4_d1 <= p3_d1;
      p4_d2 <= p3_d2;
      p4_d3 <= p3_d3;
      p4_d4 <= p3_d4;

      p5_d0 <= p4_d0;
      p5_d1 <= p4_d1;
      p5_d2 <= p4_d2;
      p5_d3 <= p4_d3;
      p5_d4 <= p4_d4;

    end

  end


  //   always @(negedge clk) begin
  //     if (s_all_en == 1) begin
  //       sum_a = sum1 + sum2 + sum3 + sum4 + sum5;
  //     end else if (accum_en == 1) begin
  //       sum_a = sum_a - sum5;
  //       sum_a = sum_a + sum1;
  //     end else begin
  //       sum_a = 0;
  //     end
  //   end

  assign sum_a = (s_all_en == 1) ? (sum1 + sum2 + sum3 +sum4 + sum5) : (accum_en == 1 ?  (sum_a - sum5 + sum1) : 0);
endmodule
