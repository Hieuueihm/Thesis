module top_module__controller (
    input clk,
    input rst_n,
    input finish_i,
    input start_i,
    input read_finish,
    output reg o_intr,
    output reg read_en
);
  parameter IDLE = 2'b00, PROCESS = 2'b01, READ = 2'b10, FIniSH = 2'b11;
  reg [1:0] current_state, next_state;

  always @(posedge clk) begin
    if (~rst_n) current_state <= IDLE;
    else current_state <= next_state;
  end
  always @(*) begin
    case (current_state)
      IDLE:    next_state = (start_i) ? PROCESS : IDLE;
      PROCESS: next_state = (finish_i) ? READ : PROCESS;
      READ:    next_state = (read_finish) ? FIniSH : READ;
      FIniSH:  next_state = IDLE;

    endcase
  end
  always @(*) begin
    case (current_state)
      IDLE: begin
        read_en <= 0;
        o_intr  <= 0;
      end
      PROCESS: begin
      end
      READ: begin
        read_en <= 1'b1;
      end

      FIniSH: begin
        read_en <= 1'b0;
        o_intr  <= 1'b1;
      end


    endcase

  end




endmodule
