module Median_filter_9x9 #(parameter ROWS = 11,
                           parameter COLS = 11)
                          (input clk,
                           input rst,
                           input done_i,
                           input [7:0] d0_i,
                           input [7:0] d1_i,
                           input [7:0] d2_i,
                           input [7:0] d3_i,
                           input [7:0] d4_i,
                           input [7:0] d5_i,
                           input [7:0] d6_i,
                           input [7:0] d7_i,
                           input [7:0] d8_i,
                           output [7:0] median_o,
                           output done_o);
    wire [7:0] data0,
    data1,
    data2,
    data3,
    data4,
    data5,
    data6,
    data7,
    data8,
    data9,
    data10,
    data11,
    data12,
    data13,
    data14,
    data15,
    data16,
    data17,
    data18,
    data19,
    data20,
    data21,
    data22,
    data23,
    data24,
    data25,
    data26,
    data27,
    data28,
    data29,
    data30,
    data31,
    data32,
    data33,
    data34,
    data35,
    data36,
    data37,
    data38,
    data39,
    data40,
    data41,
    data42,
    data43,
    data44,
    data45,
    data46,
    data47,
    data48,
    data49,
    data50,
    data51,
    data52,
    data53,
    data54,
    data55,
    data56,
    data57,
    data58,
    data59,
    data60,
    data61,
    data62,
    data63,
    data64,
    data65,
    data66,
    data67,
    data68,
    data69,
    data70,
    data71,
    data72,
    data73,
    data74,
    data75,
    data76,
    data77,
    data78,
    data79,
    data80;
    wire done_o_modulate;
    Data_modulate_9x9 #(
    .ROWS(ROWS),
    .COLS(COLS)
    ) MEDIAN_9X9_DATA_MODULATE (
    .clk(clk),
    .rst(rst),
    .d0_i(d0_i),  // 99
    .d1_i(d1_i),  // 8
    .d2_i(d2_i),  // 7
    .d3_i(d3_i),
    .d4_i(d4_i),
    .d5_i(d5_i),
    .d6_i(d6_i),
    .d7_i(d7_i),
    .d8_i(d8_i),
    // d5 d4 d3
    .done_i(done_i),
    .d0_o(data0),
    .d1_o(data1),
    .d2_o(data2),
    .d3_o(data3),
    .d4_o(data4),
    .d5_o(data5),
    .d6_o(data6),
    .d7_o(data7),
    .d8_o(data8),
    .d9_o(data9),
    .d10_o(data10),
    .d11_o(data11),
    .d12_o(data12),
    .d13_o(data13),
    .d14_o(data14),
    .d15_o(data15),
    .d16_o(data16),
    .d17_o(data17),
    .d18_o(data18),
    .d19_o(data19),
    .d20_o(data20),
    .d21_o(data21),
    .d22_o(data22),
    .d23_o(data23),
    .d24_o(data24),
    .d25_o(data25),
    .d26_o(data26),
    .d27_o(data27),
    .d28_o(data28),
    .d29_o(data29),
    .d30_o(data30),
    .d31_o(data31),
    .d32_o(data32),
    .d33_o(data33),
    .d34_o(data34),
    .d35_o(data35),
    .d36_o(data36),
    .d37_o(data37),
    .d38_o(data38),
    .d39_o(data39),
    .d40_o(data40),
    .d41_o(data41),
    .d42_o(data42),
    .d43_o(data43),
    .d44_o(data44),
    .d45_o(data45),
    .d46_o(data46),
    .d47_o(data47),
    .d48_o(data48),
    .d49_o(data49),
    .d50_o(data50),
    .d51_o(data51),
    .d52_o(data52),
    .d53_o(data53),
    .d54_o(data54),
    .d55_o(data55),
    .d56_o(data56),
    .d57_o(data57),
    .d58_o(data58),
    .d59_o(data59),
    .d60_o(data60),
    .d61_o(data61),
    .d62_o(data62),
    .d63_o(data63),
    .d64_o(data64),
    .d65_o(data65),
    .d66_o(data66),
    .d67_o(data67),
    .d68_o(data68),
    .d69_o(data69),
    .d70_o(data70),
    .d71_o(data71),
    .d72_o(data72),
    .d73_o(data73),
    .d74_o(data74),
    .d75_o(data75),
    .d76_o(data76),
    .d77_o(data77),
    .d78_o(data78),
    .d79_o(data79),
    .d80_o(data80),
    
    
    
    .done_o(done_o_modulate)
    
    );
    
    Median_filter_9x9_calc MEDIAN_9x9_CALC (
    .clk(clk),
    .rst(rst),
    .done_i(done_o_modulate),
    .S1(data0),
    .S2(data1),
    .S3(data2),
    .S4(data3),
    .S5(data4),
    .S6(data5),
    .S7(data6),
    .S8(data7),
    
    .S9 (data8),
    .S10(data9),
    .S11(data10),
    .S12(data11),
    .S13(data12),
    .S14(data13),
    .S15(data14),
    .S16(data15),
    .S17(data16),
    .S18(data17),
    .S19(data18),
    .S20(data19),
    .S21(data20),
    .S22(data21),
    .S23(data22),
    .S24(data23),
    .S25(data24),
    .S26(data25),
    .S27(data26),
    .S28(data27),
    .S29(data28),
    .S30(data29),
    .S31(data30),
    .S32(data31),
    .S33(data32),
    .S34(data33),
    .S35(data34),
    .S36(data35),
    .S37(data36),
    .S38(data37),
    .S39(data38),
    .S40(data39),
    .S41(data40),
    .S42(data41),
    .S43(data42),
    .S44(data43),
    .S45(data44),
    .S46(data45),
    .S47(data46),
    .S48(data47),
    .S49(data48),
    .S50(data49),
    .S51(data50),
    .S52(data51),
    .S53(data52),
    .S54(data53),
    .S55(data54),
    .S56(data55),
    .S57(data56),
    .S58(data57),
    .S59(data58),
    .S60(data59),
    .S61(data60),
    .S62(data61),
    .S63(data62),
    .S64(data63),
    .S65(data64),
    .S66(data65),
    .S67(data66),
    .S68(data67),
    .S69(data68),
    .S70(data69),
    .S71(data70),
    .S72(data71),
    .S73(data72),
    .S74(data73),
    .S75(data74),
    .S76(data75),
    .S77(data76),
    .S78(data77),
    .S79(data78),
    .S80(data79),
    .S81(data80),
    
    
    
    .median_o(median_o),
    .done_o  (done_o)
    );
    
    
    
endmodule
