module Window_buffer_5x5 #(parameter COLS = 7,
                           parameter ROWS = 7)
                          (input clk,
                           input rst_n,
                           input done_i,
                           input[7:0] S1_i,
                           S2_i,
                           S3_i,
                           S4_i,
                           S5_i,
                           output[7:0] S1_o,
                           S2_o,
                           S3_o,
                           S4_o,
                           S5_o,
                           S6_o,
                           S7_o,
                           S8_o,
                           S9_o,
                           S10_o,
                           S11_o,
                           S12_o,
                           S13_o,
                           S14_o,
                           S15_o,
                           S16_o,
                           S17_o,
                           S18_o,
                           S19_o,
                           S20_o,
                           S21_o,
                           S22_o,
                           S23_o,
                           S24_o,
                           S25_o,
                           output done_o,
                           output progress_done_o);
    wire i_row_eq_max, i_col_eq_max, i_col_ge_threshold;
    wire count_en;
    Window_buffer_5x5_controller WINDOW_BUFFER_5X5_CONTROLLER(
    .clk(clk),
    .rst_n(rst_n),
    .done_i(done_i),
    .i_row_eq_max(i_row_eq_max),
    .i_col_eq_max(i_col_eq_max),
    .i_col_ge_threshold(i_col_ge_threshold),
    .count_en(count_en),
    .progress_done(progress_done_o),
    .done_o(done_o));
    
    Window_buffer_5x5_datapath #(.COLS(COLS),
    .ROWS(ROWS))
    WINDOW_BUFFER_5X5_DATAPATH
    (
    .clk(clk),
    .rst_n(rst_n),
    .count_en(count_en),
    .S1_i(S1_i),
    .S2_i(S2_i),
    .S3_i(S3_i),
    .S4_i(S4_i),
    .S5_i(S5_i),
    .i_row_eq_max(i_row_eq_max),
    .S1_o(S1_o),
    .S2_o(S2_o),
    .S3_o(S3_o),
    .S4_o(S4_o),
    .S5_o(S5_o),
    .S6_o(S6_o),
    .S7_o(S7_o),
    .S8_o(S8_o),
    .S9_o(S9_o),
    .S10_o(S10_o),
    .S11_o(S11_o),
    .S12_o(S12_o),
    .S13_o(S13_o),
    .S14_o(S14_o),
    .S15_o(S15_o),
    .S16_o(S16_o),
    .S17_o(S17_o),
    .S18_o(S18_o),
    .S19_o(S19_o),
    .S20_o(S20_o),
    .S21_o(S21_o),
    .S22_o(S22_o),
    .S23_o(S23_o),
    .S24_o(S24_o),
    .S25_o(S25_o),
    .i_col_eq_max(i_col_eq_max),
    .i_col_ge_threshold(i_col_ge_threshold));
    
endmodule
